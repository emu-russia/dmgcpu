module PPU2 (  cclk, clk6, n_reset2, a, d, n_oamb, oam_bl_pch, oa, n_oam_rd, n_oamb_wr, n_oama_wr, n_oama, CONST0, n_dma_phi, 
	dma_a, dma_run, 
	soc_wr, soc_rd, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, n_ppu_hard_reset, 
	nma, fexx, ff43, ff42, sprite_x_flip, sprite_x_match, bp_sel, ppu_mode3, 
	md, oam_din, v, FF43_D1, FF43_D0, n_ppu_clk, FF43_D2, h, ppu_mode2, vbl, stop_oam_eval, obj_color, vclk2, h_restart, obj_prio_ck, obj_prio, n_ppu_reset, 
	n_vram_to_oam, n_dma_phi2_latched, FF40_D3, FF40_D2, in_window, 
	FF40_D1, dma_addr_ext, sp_bp_cys, cpu_vram_oam_rd, oam_dma_wr, clk6_delay, oam_mode3_bl_pch, bp_cy, tm_cy, oam_mode3_nrd, ma0, oam_rd_ck, oam_xattr_latch_cck, oam_addr_ck);

	input wire cclk;
	input wire clk6;
	input wire n_reset2;
	input wire [7:0] a;
	inout wire [7:0] d;
	inout wire [7:0] n_oamb;
	output wire oam_bl_pch;
	output wire [7:1] oa; 		// ⚠️ lsb=1
	output wire n_oam_rd;
	output wire n_oamb_wr;
	output wire n_oama_wr;
	inout wire [7:0] n_oama;
	inout wire CONST0;
	input wire n_dma_phi;
	input wire [12:0] dma_a;
	input wire dma_run;
	input wire soc_wr;
	input wire soc_rd;
	output wire ppu_rd;
	output wire ppu_wr;
	output wire ppu_clk;
	input wire vram_to_oam;
	output wire n_ppu_hard_reset;
	inout wire [12:0] nma;
	input wire fexx;
	input wire ff43;
	input wire ff42;
	output wire sprite_x_flip;
	output wire sprite_x_match;
	input wire bp_sel;
	input wire ppu_mode3;
	inout wire [7:0] md;
	output wire FF43_D1;
	output wire FF43_D0;
	output wire n_ppu_clk;
	output wire FF43_D2;
	output wire ppu_mode2;
	input wire vbl;
	output wire stop_oam_eval;
	output wire obj_color;
	input wire vclk2;
	output wire obj_prio;
	input wire n_ppu_reset;
	input wire FF40_D3;
	input wire FF40_D2;
	input wire in_window;
	input wire FF40_D1;
	input wire sp_bp_cys;
	input wire cpu_vram_oam_rd;
	output wire clk6_delay;
	input wire bp_cy;
	input wire tm_cy;
	input wire [7:0] oam_din;
	input wire dma_addr_ext;
	input wire oam_dma_wr;
	input wire obj_prio_ck;
	input wire n_dma_phi2_latched;
	input wire ma0;
	output wire h_restart;
	output wire n_vram_to_oam;
	input wire oam_mode3_nrd;
	input wire oam_mode3_bl_pch;
	input wire oam_rd_ck;
	input wire oam_xattr_latch_cck;
	input wire oam_addr_ck;

	// H/V
	input wire [7:0] h;
	input wire [7:0] v;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;

	assign w139 = oam_din[0];
	assign w138 = vram_to_oam;
	assign w561 = oam_din[5];
	assign ppu_clk = w391;
	assign w560 = soc_rd;
	assign w551 = dma_addr_ext;
	assign w548 = n_dma_phi;
	assign w549 = clk6;
	assign n_ppu_hard_reset = w11;
	assign w161 = n_reset2;
	assign clk6_delay = w452;
	assign w160 = soc_wr;
	assign w552 = dma_a[9];
	assign w455 = dma_run;
	assign w135 = dma_a[12];
	assign w136 = dma_a[8];
	assign w50 = dma_a[4];
	assign w51 = dma_a[11];
	assign w451 = dma_a[3];
	assign w116 = dma_a[7];
	assign w115 = cpu_vram_oam_rd;
	assign w645 = dma_a[10];
	assign w404 = dma_a[5];
	assign w233 = dma_a[1];
	assign w644 = dma_a[2];
	assign w132 = dma_a[6];
	assign w131 = a[4];
	assign w553 = a[2];
	assign w499 = a[0];
	assign w498 = a[1];
	assign w124 = oam_dma_wr;
	assign w904 = a[3];
	assign w642 = a[7];
	assign w643 = a[5];
	assign w703 = dma_a[0];
	assign w46 = a[6];
	assign w564 = cclk;
	assign d[2] = w402;
	assign d[0] = w234;
	assign d[1] = w158;
	assign d[7] = w521;
	assign d[4] = w185;
	assign d[3] = w12;
	assign d[6] = w7;
	assign d[5] = w6;
	assign oa[1] = w886;
	assign CONST0 = w69;
	assign oa[2] = w148;
	assign oa[3] = w147;
	assign n_oama[5] = w164;
	assign n_oamb_wr = w127;
	assign oa[5] = w128;
	assign oa[6] = w129;
	assign oa[4] = w130;
	assign n_oama_wr = w556;
	assign n_oama[2] = w9;
	assign n_oama[3] = w163;
	assign oa[7] = w555;
	assign n_oama[1] = w60;
	assign n_oama[6] = w465;
	assign n_oama[4] = w141;
	assign n_oam_rd = w179;
	assign n_oama[0] = w510;
	assign n_oama[7] = w59;
	assign oam_bl_pch = w58;
	assign n_oamb[3] = w243;
	assign n_oamb[4] = w178;
	assign n_oamb[5] = w5;
	assign n_oamb[1] = w460;
	assign n_oamb[6] = w567;
	assign n_oamb[2] = w63;
	assign n_oamb[0] = w169;
	assign n_oamb[7] = w168;
	assign w571 = n_ppu_reset;
	assign w200 = h[6];
	assign w199 = obj_prio_ck;
	assign h_restart = w409;
	assign stop_oam_eval = w569;
	assign obj_prio = w97;
	assign w859 = vbl;
	assign w423 = h[0];
	assign w96 = h[1];
	assign w408 = vclk2;
	assign w858 = tm_cy;
	assign w54 = FF40_D1;
	assign w55 = oam_xattr_latch_cck;
	assign w697 = h[5];
	assign w399 = h[2];
	assign w171 = ma0;
	assign obj_color = w419;
	assign w172 = oam_mode3_nrd;
	assign w914 = bp_sel;
	assign w492 = oam_addr_ck;
	assign w108 = FF40_D3;
	assign w862 = in_window;
	assign w109 = FF40_D2;
	assign FF43_D2 = w400;
	assign w188 = h[4];
	assign w389 = v[0];
	assign w439 = v[1];
	assign w230 = h[3];
	assign n_ppu_clk = w390;
	assign FF43_D0 = w422;
	assign ppu_mode2 = w3;
	assign w815 = oam_rd_ck;
	assign w155 = bp_cy;
	assign FF43_D1 = w156;
	assign sprite_x_match = w545;
	assign w546 = oam_mode3_bl_pch;
	assign w912 = sp_bp_cys;
	assign nma[2] = w52;
	assign md[6] = w458;
	assign md[0] = w143;
	assign ppu_wr = w205;
	assign md[7] = w173;
	assign sprite_x_flip = w174;
	assign md[4] = w142;
	assign md[1] = w61;
	assign nma[10] = w107;
	assign md[3] = w457;
	assign w4 = ppu_mode3;
	assign md[2] = w701;
	assign w398 = v[2];
	assign nma[11] = w394;
	assign w393 = ff42;
	assign nma[5] = w405;
	assign nma[12] = w134;
	assign w539 = v[3];
	assign nma[3] = w450;
	assign w471 = v[4];
	assign nma[4] = w694;
	assign nma[0] = w702;
	assign nma[6] = w133;
	assign w447 = v[6];
	assign nma[1] = w318;
	assign w317 = v[5];
	assign w104 = h[7];
	assign nma[7] = w117;
	assign nma[8] = w118;
	assign w105 = v[7];
	assign nma[9] = w525;
	assign w526 = oam_din[2];
	assign ppu_rd = w1;
	assign w2 = ff43;
	assign w901 = oam_din[7];
	assign md[5] = w887;
	assign w207 = n_dma_phi2_latched;
	assign w454 = fexx;
	assign w527 = oam_din[1];
	assign w534 = oam_din[4];
	assign w558 = oam_din[6];
	assign n_vram_to_oam = w559;
	assign w562 = oam_din[3];

	// Instances

	dmg_not g1 (.a(w138), .x(w559) );
	dmg_not g2 (.a(w454), .x(w456) );
	dmg_not g3 (.a(w532), .x(w443) );
	dmg_not g4 (.a(w492), .x(w459) );
	dmg_not g5 (.a(w862), .x(w857) );
	dmg_not g6 (.a(w859), .x(w407) );
	dmg_not g7 (.a(w174), .x(w433) );
	dmg_not g8 (.a(w570), .x(w712) );
	dmg_not g9 (.a(w571), .x(w570) );
	dmg_not g10 (.a(w571), .x(w688) );
	dmg_not g11 (.a(w297), .x(w295) );
	dmg_not g12 (.a(w409), .x(w410) );
	dmg_not g13 (.a(w297), .x(w717) );
	dmg_not g14 (.a(w875), .x(w722) );
	dmg_not g15 (.a(w266), .x(w875) );
	dmg_not g16 (.a(w220), .x(w270) );
	dmg_not g17 (.a(w574), .x(w221) );
	dmg_not g18 (.a(w219), .x(w218) );
	dmg_not g19 (.a(w292), .x(w293) );
	dmg_not g20 (.a(w293), .x(w40) );
	dmg_not g21 (.a(w266), .x(w265) );
	dmg_not g22 (.a(w226), .x(w227) );
	dmg_not g23 (.a(w295), .x(w296) );
	dmg_not g24 (.a(w811), .x(w184) );
	dmg_not g25 (.a(w550), .x(w452) );
	dmg_not g26 (.a(w184), .x(w10) );
	dmg_not g27 (.a(w348), .x(w489) );
	dmg_not g28 (.a(w389), .x(w388) );
	dmg_not g29 (.a(w321), .x(w320) );
	dmg_not g30 (.a(w227), .x(w747) );
	dmg_not g31 (.a(w337), .x(w372) );
	dmg_not g32 (.a(w575), .x(w300) );
	dmg_not g33 (.a(w215), .x(w824) );
	dmg_not g34 (.a(w221), .x(w272) );
	dmg_not g35 (.a(w343), .x(w341) );
	dmg_not g36 (.a(w215), .x(w214) );
	dmg_not g37 (.a(w513), .x(w292) );
	dmg_not g38 (.a(w369), .x(w512) );
	dmg_not g39 (.a(w197), .x(w39) );
	dmg_not g40 (.a(w662), .x(w664) );
	dmg_not g41 (.a(w913), .x(w666) );
	dmg_not g42 (.a(w633), .x(w753) );
	dmg_not g43 (.a(w333), .x(w334) );
	dmg_not g44 (.a(w750), .x(w766) );
	dmg_not g45 (.a(w768), .x(w803) );
	dmg_not g46 (.a(w381), .x(w802) );
	dmg_not g47 (.a(w666), .x(w432) );
	dmg_not g48 (.a(w26), .x(w386) );
	dmg_not g49 (.a(w616), .x(w349) );
	dmg_not g50 (.a(w479), .x(w869) );
	dmg_not g51 (.a(w473), .x(w474) );
	dmg_not g52 (.a(w476), .x(w475) );
	dmg_not g53 (.a(w817), .x(w816) );
	dmg_not g54 (.a(w485), .x(w484) );
	dmg_not g55 (.a(w482), .x(w483) );
	dmg_not g56 (.a(w105), .x(w106) );
	dmg_not g57 (.a(w58), .x(w242) );
	dmg_not g58 (.a(w349), .x(w690) );
	dmg_not g59 (.a(w363), .x(w362) );
	dmg_not g60 (.a(w15), .x(w590) );
	dmg_not g61 (.a(w214), .x(w276) );
	dmg_not g62 (.a(w603), .x(w595) );
	dmg_not g63 (.a(w595), .x(w600) );
	dmg_not g64 (.a(w64), .x(w65) );
	dmg_not g65 (.a(w738), .x(w294) );
	dmg_not g66 (.a(w690), .x(w736) );
	dmg_not g67 (.a(w885), .x(w325) );
	dmg_not g68 (.a(w497), .x(w886) );
	dmg_not g69 (.a(w146), .x(w147) );
	dmg_not g70 (.a(w500), .x(w148) );
	dmg_not g71 (.a(w554), .x(w555) );
	dmg_not g72 (.a(w641), .x(w128) );
	dmg_not g73 (.a(w49), .x(w130) );
	dmg_not g74 (.a(w841), .x(w842) );
	dmg_not g75 (.a(w165), .x(w841) );
	dmg_not g76 (.a(w237), .x(w120) );
	dmg_not g77 (.a(w58), .x(w237) );
	dmg_not g78 (.a(w511), .x(w431) );
	dmg_not g79 (.a(w843), .x(w415) );
	dmg_not g80 (.a(w349), .x(w350) );
	dmg_not g81 (.a(w344), .x(w583) );
	dmg_not g82 (.a(w344), .x(w282) );
	dmg_not g83 (.a(w282), .x(w283) );
	dmg_not g84 (.a(w661), .x(w603) );
	dmg_not g85 (.a(w291), .x(w288) );
	dmg_not g86 (.a(w70), .x(w82) );
	dmg_not g87 (.a(w321), .x(w591) );
	dmg_not g88 (.a(w591), .x(w77) );
	dmg_not g89 (.a(w692), .x(w593) );
	dmg_not g90 (.a(w583), .x(w585) );
	dmg_not g91 (.a(w603), .x(w662) );
	dmg_not g92 (.a(w365), .x(w822) );
	dmg_not g93 (.a(w746), .x(w821) );
	dmg_not g94 (.a(w623), .x(w622) );
	dmg_not g95 (.a(w632), .x(w786) );
	dmg_not g96 (.a(w321), .x(w529) );
	dmg_not g97 (.a(w350), .x(w414) );
	dmg_not g98 (.a(w837), .x(w351) );
	dmg_not g99 (.a(w666), .x(w667) );
	dmg_not g100 (.a(w15), .x(w258) );
	dmg_not g101 (.a(w667), .x(w866) );
	dmg_not g102 (.a(w631), .x(w630) );
	dmg_not g103 (.a(w529), .x(w247) );
	dmg_not g104 (.a(w242), .x(w314) );
	dmg_not g105 (.a(w508), .x(w463) );
	dmg_not g106 (.a(w447), .x(w446) );
	dmg_not g107 (.a(w471), .x(w472) );
	dmg_not g108 (.a(w317), .x(w316) );
	dmg_not g109 (.a(w539), .x(w540) );
	dmg_not g110 (.a(w349), .x(w348) );
	dmg_not g111 (.a(w398), .x(w397) );
	dmg_not g112 (.a(w109), .x(w818) );
	dmg_not g113 (.a(w292), .x(w291) );
	dmg_not g114 (.a(w666), .x(w306) );
	dmg_not g115 (.a(w215), .x(w369) );
	dmg_not g116 (.a(w306), .x(w305) );
	dmg_not g117 (.a(w300), .x(w515) );
	dmg_not g118 (.a(w270), .x(w301) );
	dmg_not g119 (.a(w344), .x(w343) );
	dmg_not g120 (.a(w345), .x(w344) );
	dmg_not g121 (.a(w824), .x(w825) );
	dmg_not g122 (.a(w302), .x(w656) );
	dmg_not g123 (.a(w226), .x(w302) );
	dmg_not g124 (.a(w216), .x(w215) );
	dmg_not g125 (.a(w322), .x(w321) );
	dmg_not g126 (.a(w265), .x(w90) );
	dmg_not g127 (.a(w22), .x(w21) );
	dmg_not g128 (.a(w757), .x(w584) );
	dmg_not g129 (.a(w371), .x(w27) );
	dmg_not g130 (.a(w894), .x(w787) );
	dmg_not g131 (.a(w432), .x(w437) );
	dmg_not g132 (.a(w438), .x(w311) );
	dmg_not g133 (.a(w439), .x(w312) );
	dmg_not g134 (.a(w543), .x(w544) );
	dmg_not g135 (.a(w68), .x(w67) );
	dmg_not g136 (.a(w161), .x(w162) );
	dmg_not g137 (.a(w549), .x(w550) );
	dmg_not g138 (.a(w452), .x(w453) );
	dmg_not g139 (.a(w455), .x(w101) );
	dmg_not g140 (.a(w443), .x(w159) );
	dmg_not g141 (.a(w102), .x(w444) );
	dmg_not g142 (.a(w204), .x(w203) );
	dmg_not g143 (.a(w144), .x(w145) );
	dmg_not g144 (.a(w166), .x(w165) );
	dmg_not g145 (.a(w320), .x(w251) );
	dmg_not g146 (.a(w154), .x(w153) );
	dmg_not g147 (.a(w209), .x(w208) );
	dmg_not g148 (.a(w253), .x(w252) );
	dmg_not g149 (.a(w650), .x(w253) );
	dmg_not g150 (.a(w97), .x(w594) );
	dmg_not g151 (.a(w687), .x(w371) );
	dmg_not g152 (.a(w324), .x(w685) );
	dmg_not g153 (.a(w292), .x(w324) );
	dmg_not g154 (.a(w297), .x(w725) );
	dmg_not g155 (.a(w298), .x(w297) );
	dmg_not g156 (.a(w725), .x(w728) );
	dmg_not g157 (.a(w717), .x(w715) );
	dmg_not g158 (.a(w830), .x(w328) );
	dmg_not g159 (.a(w266), .x(w830) );
	dmg_not g160 (.a(w267), .x(w266) );
	dmg_not g161 (.a(w579), .x(w578) );
	dmg_not g162 (.a(w226), .x(w579) );
	dmg_latchnq_comp g163 (.n_ena(w579), .d(w310), .ena(w578), .nq(w827) );
	dmg_latchnq_comp g164 (.n_ena(w579), .d(w259), .ena(w578), .nq(w828) );
	dmg_latchnq_comp g165 (.n_ena(w579), .d(w66), .ena(w578), .nq(w580) );
	dmg_latchnq_comp g166 (.n_ena(w579), .d(w257), .ena(w578), .nq(w577) );
	dmg_latchnq_comp g167 (.n_ena(w830), .d(w259), .ena(w328), .nq(w327) );
	dmg_latchnq_comp g168 (.n_ena(w830), .d(w66), .ena(w328), .nq(w831) );
	dmg_latchnq_comp g169 (.n_ena(w830), .d(w257), .ena(w328), .nq(w832) );
	dmg_latchnq_comp g170 (.n_ena(w830), .d(w310), .ena(w328), .nq(w329) );
	dmg_latchnq_comp g171 (.n_ena(w717), .d(w257), .ena(w715), .nq(w720) );
	dmg_latchnq_comp g172 (.n_ena(w717), .d(w66), .ena(w715), .nq(w718) );
	dmg_latchnq_comp g173 (.n_ena(w717), .d(w310), .ena(w715), .nq(w719) );
	dmg_latchnq_comp g174 (.n_ena(w717), .d(w259), .ena(w715), .nq(w716) );
	dmg_latchnq_comp g175 (.n_ena(w875), .d(w323), .ena(w722), .nq(w878) );
	dmg_latchnq_comp g176 (.n_ena(w875), .d(w347), .ena(w722), .nq(w879) );
	dmg_latchnq_comp g177 (.n_ena(w343), .d(w66), .ena(w341), .nq(w581) );
	dmg_latchnq_comp g178 (.n_ena(w824), .d(w259), .ena(w825), .nq(w273) );
	dmg_latchnq_comp g179 (.n_ena(w725), .d(w213), .ena(w728), .nq(w880) );
	dmg_latchnq_comp g180 (.n_ena(w725), .d(w487), .ena(w728), .nq(w726) );
	dmg_latchnq_comp g181 (.n_ena(w725), .d(w347), .ena(w728), .nq(w727) );
	dmg_latchnq_comp g182 (.n_ena(w725), .d(w323), .ena(w728), .nq(w874) );
	dmg_latchnq_comp g183 (.n_ena(w725), .d(w279), .ena(w728), .nq(w873) );
	dmg_latchnq_comp g184 (.n_ena(w725), .d(w284), .ena(w728), .nq(w895) );
	dmg_latchnq_comp g185 (.n_ena(w320), .d(w257), .ena(w251), .nq(w256) );
	dmg_latchnq_comp g186 (.n_ena(w320), .d(w259), .ena(w251), .nq(w700) );
	dmg_latchnq_comp g187 (.n_ena(w320), .d(w310), .ena(w251), .nq(w853) );
	dmg_latchnq_comp g188 (.n_ena(w320), .d(w66), .ena(w251), .nq(w250) );
	dmg_latchnq_comp g189 (.n_ena(w302), .d(w284), .ena(w656), .nq(w681) );
	dmg_latchnq_comp g190 (.n_ena(w302), .d(w279), .ena(w656), .nq(w682) );
	dmg_latchnq_comp g191 (.n_ena(w302), .d(w323), .ena(w656), .nq(w683) );
	dmg_latchnq_comp g192 (.n_ena(w302), .d(w487), .ena(w656), .nq(w684) );
	dmg_latchnq_comp g193 (.n_ena(w302), .d(w347), .ena(w656), .nq(w826) );
	dmg_latchnq_comp g194 (.n_ena(w824), .d(w257), .ena(w825), .nq(w658) );
	dmg_latchnq_comp g195 (.n_ena(w302), .d(w213), .ena(w656), .nq(w657) );
	dmg_latchnq_comp g196 (.n_ena(w306), .d(w279), .ena(w305), .nq(w303) );
	dmg_latchnq_comp g197 (.n_ena(w306), .d(w284), .ena(w305), .nq(w309) );
	dmg_latchnq_comp g198 (.n_ena(w306), .d(w487), .ena(w305), .nq(w870) );
	dmg_latchnq_comp g199 (.n_ena(w662), .d(w347), .ena(w664), .nq(w691) );
	dmg_latchnq_comp g200 (.n_ena(w662), .d(w323), .ena(w664), .nq(w769) );
	dmg_latchnq_comp g201 (.n_ena(w662), .d(w284), .ena(w664), .nq(w819) );
	dmg_latchnq_comp g202 (.n_ena(w662), .d(w487), .ena(w664), .nq(w823) );
	dmg_latchnq_comp g203 (.n_ena(w242), .d(w420), .ena(w314), .nq(w419) );
	dmg_latchnq_comp g204 (.n_ena(w237), .d(w240), .ena(w120), .nq(w445) );
	dmg_latchnq_comp g205 (.n_ena(w237), .d(w111), .ena(w120), .nq(w110) );
	dmg_latchnq_comp g206 (.n_ena(w237), .d(w236), .ena(w120), .nq(w387) );
	dmg_latchnq_comp g207 (.n_ena(w237), .d(w461), .ena(w120), .nq(w313) );
	dmg_latchnq_comp g208 (.n_ena(w529), .d(w347), .ena(w247), .nq(w248) );
	dmg_latchnq_comp g209 (.n_ena(w529), .d(w487), .ena(w247), .nq(w865) );
	dmg_latchnq_comp g210 (.n_ena(w529), .d(w323), .ena(w247), .nq(w530) );
	dmg_latchnq_comp g211 (.n_ena(w529), .d(w284), .ena(w247), .nq(w838) );
	dmg_latchnq_comp g212 (.n_ena(w529), .d(w279), .ena(w247), .nq(w839) );
	dmg_latchnq_comp g213 (.n_ena(w667), .d(w66), .ena(w866), .nq(w868) );
	dmg_latchnq_comp g214 (.n_ena(w667), .d(w257), .ena(w866), .nq(w867) );
	dmg_latchnq_comp g215 (.n_ena(w667), .d(w310), .ena(w866), .nq(w733) );
	dmg_latchnq_comp g216 (.n_ena(w291), .d(w259), .ena(w288), .nq(w770) );
	dmg_latchnq_comp g217 (.n_ena(w291), .d(w310), .ena(w288), .nq(w772) );
	dmg_latchnq_comp g218 (.n_ena(w282), .d(w279), .ena(w283), .nq(w287) );
	dmg_latchnq_comp g219 (.n_ena(w282), .d(w213), .ena(w283), .nq(w281) );
	dmg_latchnq_comp g220 (.n_ena(w282), .d(w323), .ena(w283), .nq(w655) );
	dmg_latchnq_comp g221 (.n_ena(w282), .d(w347), .ena(w283), .nq(w653) );
	dmg_latchnq_comp g222 (.n_ena(w214), .d(w284), .ena(w276), .nq(w285) );
	dmg_latchnq_comp g223 (.n_ena(w64), .d(w257), .ena(w65), .nq(w739) );
	dmg_latchnq_comp g224 (.n_ena(w64), .d(w259), .ena(w65), .nq(w244) );
	dmg_latchnq_comp g225 (.n_ena(w64), .d(w310), .ena(w65), .nq(w776) );
	dmg_latchnq_comp g226 (.n_ena(w64), .d(w66), .ena(w65), .nq(w844) );
	dmg_latchnq_comp g227 (.n_ena(w690), .d(w257), .ena(w736), .nq(w735) );
	dmg_latchnq_comp g228 (.n_ena(w690), .d(w310), .ena(w736), .nq(w734) );
	dmg_latchnq_comp g229 (.n_ena(w690), .d(w259), .ena(w736), .nq(w737) );
	dmg_latchnq_comp g230 (.n_ena(w690), .d(w66), .ena(w736), .nq(w326) );
	dmg_latchnq_comp g231 (.n_ena(w242), .d(w506), .ena(w314), .nq(w511) );
	dmg_latchnq_comp g232 (.n_ena(w242), .d(w501), .ena(w314), .nq(w885) );
	dmg_latchnq_comp g233 (.n_ena(w242), .d(w502), .ena(w314), .nq(w843) );
	dmg_latchnq_comp g234 (.n_ena(w237), .d(w705), .ena(w120), .nq(w395) );
	dmg_latchnq_comp g235 (.n_ena(w237), .d(w121), .ena(w120), .nq(w396) );
	dmg_latchnq_comp g236 (.n_ena(w237), .d(w566), .ena(w120), .nq(w119) );
	dmg_latchnq_comp g237 (.n_ena(w242), .d(w14), .ena(w314), .nq(w15) );
	dmg_latchnq_comp g238 (.n_ena(w242), .d(w505), .ena(w314), .nq(w738) );
	dmg_latchnq_comp g239 (.n_ena(w667), .d(w259), .ena(w866), .nq(w668) );
	dmg_latchnq_comp g240 (.n_ena(w291), .d(w257), .ena(w288), .nq(w289) );
	dmg_latchnq_comp g241 (.n_ena(w291), .d(w66), .ena(w288), .nq(w589) );
	dmg_latchnq_comp g242 (.n_ena(w214), .d(w279), .ena(w276), .nq(w275) );
	dmg_latchnq_comp g243 (.n_ena(w282), .d(w284), .ena(w283), .nq(w286) );
	dmg_latchnq_comp g244 (.n_ena(w214), .d(w487), .ena(w276), .nq(w892) );
	dmg_latchnq_comp g245 (.n_ena(w214), .d(w323), .ena(w276), .nq(w891) );
	dmg_latchnq_comp g246 (.n_ena(w282), .d(w487), .ena(w283), .nq(w654) );
	dmg_latchnq_comp g247 (.n_ena(w214), .d(w277), .ena(w276), .nq(w278) );
	dmg_latchnq_comp g248 (.n_ena(w214), .d(w213), .ena(w276), .nq(w659) );
	dmg_latchnq_comp g249 (.n_ena(w529), .d(w213), .ena(w247), .nq(w246) );
	dmg_latchnq_comp g250 (.n_ena(w237), .d(w241), .ena(w120), .nq(w315) );
	dmg_latchnq_comp g251 (.n_ena(w662), .d(w213), .ena(w664), .nq(w85) );
	dmg_latchnq_comp g252 (.n_ena(w662), .d(w279), .ena(w664), .nq(w663) );
	dmg_latchnq_comp g253 (.n_ena(w306), .d(w323), .ena(w305), .nq(w308) );
	dmg_latchnq_comp g254 (.n_ena(w306), .d(w213), .ena(w305), .nq(w307) );
	dmg_latchnq_comp g255 (.n_ena(w306), .d(w347), .ena(w305), .nq(w680) );
	dmg_latchnq_comp g256 (.n_ena(w824), .d(w66), .ena(w825), .nq(w582) );
	dmg_latchnq_comp g257 (.n_ena(w343), .d(w259), .ena(w341), .nq(w871) );
	dmg_latchnq_comp g258 (.n_ena(w343), .d(w310), .ena(w341), .nq(w340) );
	dmg_latchnq_comp g259 (.n_ena(w343), .d(w257), .ena(w341), .nq(w342) );
	dmg_latchnq_comp g260 (.n_ena(w348), .d(w279), .ena(w489), .nq(w849) );
	dmg_latchnq_comp g261 (.n_ena(w348), .d(w323), .ena(w489), .nq(w850) );
	dmg_latchnq_comp g262 (.n_ena(w348), .d(w213), .ena(w489), .nq(w851) );
	dmg_latchnq_comp g263 (.n_ena(w242), .d(w905), .ena(w314), .nq(w97) );
	dmg_latchnq_comp g264 (.n_ena(w348), .d(w487), .ena(w489), .nq(w906) );
	dmg_latchnq_comp g265 (.n_ena(w348), .d(w347), .ena(w489), .nq(w488) );
	dmg_latchnq_comp g266 (.n_ena(w348), .d(w284), .ena(w489), .nq(w636) );
	dmg_latchnq_comp g267 (.n_ena(w242), .d(w175), .ena(w314), .nq(w174) );
	dmg_latchnq_comp g268 (.n_ena(w324), .d(w279), .ena(w685), .nq(w899) );
	dmg_latchnq_comp g269 (.n_ena(w324), .d(w347), .ena(w685), .nq(w900) );
	dmg_latchnq_comp g270 (.n_ena(w324), .d(w487), .ena(w685), .nq(w896) );
	dmg_latchnq_comp g271 (.n_ena(w324), .d(w323), .ena(w685), .nq(w686) );
	dmg_latchnq_comp g272 (.n_ena(w324), .d(w213), .ena(w685), .nq(w729) );
	dmg_latchnq_comp g273 (.n_ena(w324), .d(w284), .ena(w685), .nq(w724) );
	dmg_latchnq_comp g274 (.n_ena(w875), .d(w279), .ena(w722), .nq(w723) );
	dmg_latchnq_comp g275 (.n_ena(w875), .d(w213), .ena(w722), .nq(w876) );
	dmg_latchnq_comp g276 (.n_ena(w875), .d(w284), .ena(w722), .nq(w877) );
	dmg_latchnq_comp g277 (.n_ena(w875), .d(w487), .ena(w722), .nq(w721) );
	dmg_latchnq_comp g278 (.n_ena(w824), .d(w310), .ena(w825), .nq(w829) );
	dmg_notif0 g279 (.n_ena(w576), .a(w577), .x(w257) );
	dmg_notif0 g280 (.n_ena(w274), .a(w829), .x(w310) );
	dmg_notif0 g281 (.n_ena(w330), .a(w329), .x(w310) );
	dmg_notif0 g282 (.n_ena(w330), .a(w721), .x(w487) );
	dmg_notif0 g283 (.n_ena(w28), .a(w716), .x(w259) );
	dmg_notif0 g284 (.n_ena(w330), .a(w878), .x(w323) );
	dmg_notif0 g285 (.n_ena(w330), .a(w877), .x(w284) );
	dmg_notif0 g286 (.n_ena(w330), .a(w879), .x(w347) );
	dmg_notif0 g287 (.n_ena(w330), .a(w876), .x(w213) );
	dmg_notif0 g288 (.n_ena(w330), .a(w723), .x(w279) );
	dmg_notif0 g289 (.n_ena(w290), .a(w724), .x(w284) );
	dmg_notif0 g290 (.n_ena(w290), .a(w729), .x(w213) );
	dmg_notif0 g291 (.n_ena(w290), .a(w686), .x(w323) );
	dmg_notif0 g292 (.n_ena(w170), .a(w171), .x(w702) );
	dmg_notif0 g293 (.n_ena(w153), .a(w914), .x(w702) );
	dmg_notif0 g294 (.n_ena(w183), .a(w108), .x(w107) );
	dmg_notif0 g295 (.n_ena(w170), .a(w911), .x(w450) );
	dmg_notif0 g296 (.n_ena(w62), .a(w173), .x(w168) );
	dmg_notif0 g297 (.n_ena(w62), .a(w701), .x(w63) );
	dmg_notif0 g298 (.n_ena(w62), .a(w61), .x(w460) );
	dmg_notif0 g299 (.n_ena(w62), .a(w142), .x(w178) );
	dmg_notif0 g300 (.n_ena(w62), .a(w173), .x(w59) );
	dmg_notif0 g301 (.n_ena(w62), .a(w142), .x(w141) );
	dmg_notif0 g302 (.n_ena(w62), .a(w61), .x(w60) );
	dmg_notif0 g303 (.n_ena(w62), .a(w701), .x(w9) );
	dmg_notif0 g304 (.n_ena(w183), .a(w698), .x(w702) );
	dmg_notif0 g305 (.n_ena(w183), .a(w814), .x(w52) );
	dmg_notif0 g306 (.n_ena(w183), .a(w448), .x(w318) );
	dmg_notif0 g307 (.n_ena(w183), .a(w533), .x(w694) );
	dmg_notif0 g308 (.n_ena(w62), .a(w887), .x(w5) );
	dmg_notif0 g309 (.n_ena(w62), .a(w887), .x(w164) );
	dmg_notif0 g310 (.n_ena(w140), .a(w562), .x(w163) );
	dmg_notif0 g311 (.n_ena(w140), .a(w562), .x(w243) );
	dmg_notif0 g312 (.n_ena(w203), .a(w442), .x(w6) );
	dmg_notif0 g313 (.n_ena(w203), .a(w186), .x(w185) );
	dmg_notif0 g314 (.n_ena(w203), .a(w890), .x(w521) );
	dmg_notif0 g315 (.n_ena(w203), .a(w401), .x(w402) );
	dmg_notif0 g316 (.n_ena(w145), .a(w469), .x(w185) );
	dmg_notif0 g317 (.n_ena(w183), .a(w524), .x(w117) );
	dmg_notif0 g318 (.n_ena(w183), .a(w180), .x(w118) );
	dmg_notif0 g319 (.n_ena(w183), .a(w468), .x(w133) );
	dmg_notif0 g320 (.n_ena(w183), .a(w812), .x(w450) );
	dmg_notif0 g321 (.n_ena(w183), .a(w149), .x(w134) );
	dmg_notif0 g322 (.n_ena(w183), .a(w149), .x(w394) );
	dmg_notif0 g323 (.n_ena(w62), .a(w457), .x(w163) );
	dmg_notif0 g324 (.n_ena(w62), .a(w458), .x(w465) );
	dmg_notif0 g325 (.n_ena(w62), .a(w457), .x(w243) );
	dmg_notif0 g326 (.n_ena(w545), .a(w67), .x(w66) );
	dmg_notif0 g327 (.n_ena(w545), .a(w544), .x(w259) );
	dmg_notif0 g328 (.n_ena(w545), .a(w311), .x(w310) );
	dmg_notif0 g329 (.n_ena(w290), .a(w899), .x(w279) );
	dmg_notif0 g330 (.n_ena(w290), .a(w900), .x(w347) );
	dmg_notif0 g331 (.n_ena(w290), .a(w896), .x(w487) );
	dmg_notif0 g332 (.n_ena(w28), .a(w895), .x(w284) );
	dmg_notif0 g333 (.n_ena(w28), .a(w873), .x(w279) );
	dmg_notif0 g334 (.n_ena(w28), .a(w726), .x(w487) );
	dmg_notif0 g335 (.n_ena(w28), .a(w880), .x(w213) );
	dmg_notif0 g336 (.n_ena(w280), .a(w342), .x(w257) );
	dmg_notif0 g337 (.n_ena(w280), .a(w340), .x(w310) );
	dmg_notif0 g338 (.n_ena(w304), .a(w680), .x(w347) );
	dmg_notif0 g339 (.n_ena(w304), .a(w307), .x(w213) );
	dmg_notif0 g340 (.n_ena(w304), .a(w308), .x(w323) );
	dmg_notif0 g341 (.n_ena(w245), .a(w663), .x(w279) );
	dmg_notif0 g342 (.n_ena(w245), .a(w85), .x(w213) );
	dmg_notif0 g343 (.n_ena(w635), .a(w906), .x(w487) );
	dmg_notif0 g344 (.n_ena(w153), .a(w808), .x(w318) );
	dmg_notif0 g345 (.n_ena(w137), .a(w703), .x(w702) );
	dmg_notif0 g346 (.n_ena(w137), .a(w132), .x(w133) );
	dmg_notif0 g347 (.n_ena(w137), .a(w233), .x(w318) );
	dmg_notif0 g348 (.n_ena(w203), .a(w864), .x(w234) );
	dmg_notif0 g349 (.n_ena(w203), .a(w157), .x(w158) );
	dmg_notif0 g350 (.n_ena(w137), .a(w645), .x(w107) );
	dmg_notif0 g351 (.n_ena(w137), .a(w116), .x(w117) );
	dmg_notif0 g352 (.n_ena(w403), .a(w404), .x(w641) );
	dmg_notif0 g353 (.n_ena(w403), .a(w50), .x(w49) );
	dmg_notif0 g354 (.n_ena(w137), .a(w136), .x(w118) );
	dmg_notif0 g355 (.n_ena(w137), .a(w135), .x(w134) );
	dmg_notif0 g356 (.n_ena(w48), .a(w643), .x(w641) );
	dmg_notif0 g357 (.n_ena(w48), .a(w553), .x(w500) );
	dmg_notif0 g358 (.n_ena(w48), .a(w499), .x(w464) );
	dmg_notif0 g359 (.n_ena(w518), .a(w69), .x(w464) );
	dmg_notif0 g360 (.n_ena(w518), .a(w516), .x(w146) );
	dmg_notif0 g361 (.n_ena(w475), .a(w149), .x(w863) );
	dmg_notif0 g362 (.n_ena(w475), .a(w284), .x(w146) );
	dmg_notif0 g363 (.n_ena(w145), .a(w528), .x(w7) );
	dmg_notif0 g364 (.n_ena(w145), .a(w520), .x(w521) );
	dmg_notif0 g365 (.n_ena(w145), .a(w537), .x(w12) );
	dmg_notif0 g366 (.n_ena(w145), .a(w536), .x(w6) );
	dmg_notif0 g367 (.n_ena(w145), .a(w441), .x(w402) );
	dmg_notif0 g368 (.n_ena(w518), .a(w517), .x(w500) );
	dmg_notif0 g369 (.n_ena(w145), .a(w646), .x(w158) );
	dmg_notif0 g370 (.n_ena(w475), .a(w487), .x(w500) );
	dmg_notif0 g371 (.n_ena(w518), .a(w708), .x(w554) );
	dmg_notif0 g372 (.n_ena(w170), .a(w445), .x(w107) );
	dmg_notif0 g373 (.n_ena(w518), .a(w709), .x(w47) );
	dmg_notif0 g374 (.n_ena(w170), .a(w315), .x(w525) );
	dmg_notif0 g375 (.n_ena(w274), .a(w582), .x(w66) );
	dmg_notif0 g376 (.n_ena(w280), .a(w871), .x(w259) );
	dmg_notif0 g377 (.n_ena(w280), .a(w653), .x(w347) );
	dmg_notif0 g378 (.n_ena(w249), .a(w248), .x(w347) );
	dmg_notif0 g379 (.n_ena(w170), .a(w395), .x(w394) );
	dmg_notif0 g380 (.n_ena(w123), .a(w7), .x(w567) );
	dmg_notif0 g381 (.n_ena(w123), .a(w6), .x(w5) );
	dmg_notif0 g382 (.n_ena(w123), .a(w12), .x(w163) );
	dmg_notif0 g383 (.n_ena(w123), .a(w6), .x(w164) );
	dmg_notif0 g384 (.n_ena(w123), .a(w12), .x(w243) );
	dmg_notif0 g385 (.n_ena(w123), .a(w185), .x(w178) );
	dmg_notif0 g386 (.n_ena(w123), .a(w234), .x(w510) );
	dmg_notif0 g387 (.n_ena(w123), .a(w234), .x(w169) );
	dmg_notif0 g388 (.n_ena(w123), .a(w185), .x(w141) );
	dmg_notif0 g389 (.n_ena(w123), .a(w158), .x(w60) );
	dmg_notif0 g390 (.n_ena(w123), .a(w521), .x(w59) );
	dmg_notif0 g391 (.n_ena(w123), .a(w521), .x(w168) );
	dmg_notif0 g392 (.n_ena(w123), .a(w158), .x(w460) );
	dmg_notif0 g393 (.n_ena(w211), .a(w212), .x(w213) );
	dmg_notif0 g394 (.n_ena(w635), .a(w326), .x(w66) );
	dmg_notif0 g395 (.n_ena(w635), .a(w735), .x(w257) );
	dmg_notif0 g396 (.n_ena(w245), .a(w776), .x(w310) );
	dmg_notif0 g397 (.n_ena(w245), .a(w739), .x(w257) );
	dmg_notif0 g398 (.n_ena(w290), .a(w589), .x(w66) );
	dmg_notif0 g399 (.n_ena(w290), .a(w289), .x(w257) );
	dmg_notif0 g400 (.n_ena(w274), .a(w275), .x(w279) );
	dmg_notif0 g401 (.n_ena(w280), .a(w286), .x(w284) );
	dmg_notif0 g402 (.n_ena(w274), .a(w285), .x(w284) );
	dmg_notif0 g403 (.n_ena(w274), .a(w891), .x(w323) );
	dmg_notif0 g404 (.n_ena(w274), .a(w892), .x(w487) );
	dmg_notif0 g405 (.n_ena(w280), .a(w654), .x(w487) );
	dmg_notif0 g406 (.n_ena(w274), .a(w278), .x(w277) );
	dmg_notif0 g407 (.n_ena(w280), .a(w655), .x(w323) );
	dmg_notif0 g408 (.n_ena(w280), .a(w287), .x(w279) );
	dmg_notif0 g409 (.n_ena(w280), .a(w281), .x(w213) );
	dmg_notif0 g410 (.n_ena(w245), .a(w244), .x(w259) );
	dmg_notif0 g411 (.n_ena(w245), .a(w844), .x(w66) );
	dmg_notif0 g412 (.n_ena(w304), .a(w668), .x(w259) );
	dmg_notif0 g413 (.n_ena(w635), .a(w734), .x(w310) );
	dmg_notif0 g414 (.n_ena(w635), .a(w737), .x(w259) );
	dmg_notif0 g415 (.n_ena(w123), .a(w7), .x(w465) );
	dmg_notif0 g416 (.n_ena(w48), .a(w498), .x(w497) );
	dmg_notif0 g417 (.n_ena(w48), .a(w46), .x(w47) );
	dmg_notif0 g418 (.n_ena(w48), .a(w904), .x(w146) );
	dmg_notif0 g419 (.n_ena(w518), .a(w69), .x(w497) );
	dmg_notif0 g420 (.n_ena(w203), .a(w232), .x(w12) );
	dmg_notif0 g421 (.n_ena(w475), .a(w149), .x(w497) );
	dmg_notif0 g422 (.n_ena(w140), .a(w139), .x(w510) );
	dmg_notif0 g423 (.n_ena(w140), .a(w139), .x(w169) );
	dmg_notif0 g424 (.n_ena(w145), .a(w638), .x(w234) );
	dmg_notif0 g425 (.n_ena(w123), .a(w402), .x(w9) );
	dmg_notif0 g426 (.n_ena(w123), .a(w402), .x(w63) );
	dmg_notif0 g427 (.n_ena(w211), .a(w840), .x(w284) );
	dmg_notif0 g428 (.n_ena(w211), .a(w649), .x(w487) );
	dmg_notif0 g429 (.n_ena(w211), .a(w652), .x(w347) );
	dmg_notif0 g430 (.n_ena(w211), .a(w490), .x(w279) );
	dmg_notif0 g431 (.n_ena(w211), .a(w531), .x(w323) );
	dmg_notif0 g432 (.n_ena(w62), .a(w143), .x(w510) );
	dmg_notif0 g433 (.n_ena(w170), .a(w119), .x(w118) );
	dmg_notif0 g434 (.n_ena(w62), .a(w143), .x(w169) );
	dmg_notif0 g435 (.n_ena(w170), .a(w110), .x(w117) );
	dmg_notif0 g436 (.n_ena(w249), .a(w865), .x(w487) );
	dmg_notif0 g437 (.n_ena(w249), .a(w246), .x(w213) );
	dmg_notif0 g438 (.n_ena(w249), .a(w530), .x(w323) );
	dmg_notif0 g439 (.n_ena(w249), .a(w838), .x(w284) );
	dmg_notif0 g440 (.n_ena(w249), .a(w839), .x(w279) );
	dmg_notif0 g441 (.n_ena(w545), .a(w869), .x(w257) );
	dmg_notif0 g442 (.n_ena(w304), .a(w868), .x(w66) );
	dmg_notif0 g443 (.n_ena(w304), .a(w867), .x(w257) );
	dmg_notif0 g444 (.n_ena(w245), .a(w823), .x(w487) );
	dmg_notif0 g445 (.n_ena(w245), .a(w819), .x(w284) );
	dmg_notif0 g446 (.n_ena(w245), .a(w691), .x(w347) );
	dmg_notif0 g447 (.n_ena(w245), .a(w769), .x(w323) );
	dmg_notif0 g448 (.n_ena(w304), .a(w733), .x(w310) );
	dmg_notif0 g449 (.n_ena(w290), .a(w770), .x(w259) );
	dmg_notif0 g450 (.n_ena(w304), .a(w870), .x(w487) );
	dmg_notif0 g451 (.n_ena(w304), .a(w309), .x(w284) );
	dmg_notif0 g452 (.n_ena(w290), .a(w772), .x(w310) );
	dmg_notif0 g453 (.n_ena(w304), .a(w303), .x(w279) );
	dmg_notif0 g454 (.n_ena(w576), .a(w657), .x(w213) );
	dmg_notif0 g455 (.n_ena(w274), .a(w658), .x(w257) );
	dmg_notif0 g456 (.n_ena(w274), .a(w659), .x(w213) );
	dmg_notif0 g457 (.n_ena(w170), .a(w695), .x(w694) );
	dmg_notif0 g458 (.n_ena(w170), .a(w313), .x(w405) );
	dmg_notif0 g459 (.n_ena(w444), .a(w323), .x(w554) );
	dmg_notif0 g460 (.n_ena(w444), .a(w279), .x(w47) );
	dmg_notif0 g461 (.n_ena(w444), .a(w213), .x(w49) );
	dmg_notif0 g462 (.n_ena(w444), .a(w347), .x(w641) );
	dmg_notif0 g463 (.n_ena(w518), .a(w640), .x(w641) );
	dmg_notif0 g464 (.n_ena(w518), .a(w494), .x(w49) );
	dmg_notif0 g465 (.n_ena(w137), .a(w51), .x(w394) );
	dmg_notif0 g466 (.n_ena(w137), .a(w644), .x(w52) );
	dmg_notif0 g467 (.n_ena(w137), .a(w451), .x(w450) );
	dmg_notif0 g468 (.n_ena(w403), .a(w233), .x(w497) );
	dmg_notif0 g469 (.n_ena(w403), .a(w703), .x(w863) );
	dmg_notif0 g470 (.n_ena(w403), .a(w132), .x(w47) );
	dmg_notif0 g471 (.n_ena(w403), .a(w644), .x(w500) );
	dmg_notif0 g472 (.n_ena(w403), .a(w451), .x(w146) );
	dmg_notif0 g473 (.n_ena(w403), .a(w116), .x(w554) );
	dmg_notif0 g474 (.n_ena(w48), .a(w642), .x(w554) );
	dmg_notif0 g475 (.n_ena(w48), .a(w131), .x(w49) );
	dmg_notif0 g476 (.n_ena(w137), .a(w552), .x(w525) );
	dmg_notif0 g477 (.n_ena(w137), .a(w50), .x(w694) );
	dmg_notif0 g478 (.n_ena(w137), .a(w404), .x(w405) );
	dmg_notif0 g479 (.n_ena(w203), .a(w202), .x(w7) );
	dmg_notif0 g480 (.n_ena(w183), .a(w182), .x(w525) );
	dmg_notif0 g481 (.n_ena(w183), .a(w467), .x(w405) );
	dmg_notif0 g482 (.n_ena(w153), .a(w150), .x(w450) );
	dmg_notif0 g483 (.n_ena(w170), .a(w69), .x(w134) );
	dmg_notif0 g484 (.n_ena(w153), .a(w152), .x(w52) );
	dmg_notif0 g485 (.n_ena(w635), .a(w636), .x(w284) );
	dmg_notif0 g486 (.n_ena(w635), .a(w488), .x(w347) );
	dmg_notif0 g487 (.n_ena(w635), .a(w851), .x(w213) );
	dmg_notif0 g488 (.n_ena(w635), .a(w850), .x(w323) );
	dmg_notif0 g489 (.n_ena(w576), .a(w681), .x(w284) );
	dmg_notif0 g490 (.n_ena(w576), .a(w682), .x(w279) );
	dmg_notif0 g491 (.n_ena(w576), .a(w683), .x(w323) );
	dmg_notif0 g492 (.n_ena(w576), .a(w684), .x(w487) );
	dmg_notif0 g493 (.n_ena(w576), .a(w826), .x(w347) );
	dmg_notif0 g494 (.n_ena(w576), .a(w827), .x(w310) );
	dmg_notif0 g495 (.n_ena(w576), .a(w828), .x(w259) );
	dmg_notif0 g496 (.n_ena(w280), .a(w581), .x(w66) );
	dmg_notif0 g497 (.n_ena(w576), .a(w580), .x(w66) );
	dmg_notif0 g498 (.n_ena(w274), .a(w273), .x(w259) );
	dmg_notif0 g499 (.n_ena(w330), .a(w327), .x(w259) );
	dmg_notif0 g500 (.n_ena(w330), .a(w831), .x(w66) );
	dmg_notif0 g501 (.n_ena(w330), .a(w832), .x(w257) );
	dmg_notif0 g502 (.n_ena(w28), .a(w718), .x(w66) );
	dmg_notif0 g503 (.n_ena(w28), .a(w719), .x(w310) );
	dmg_notif0 g504 (.n_ena(w28), .a(w720), .x(w257) );
	dmg_notif0 g505 (.n_ena(w28), .a(w727), .x(w347) );
	dmg_notif0 g506 (.n_ena(w28), .a(w874), .x(w323) );
	dmg_notif0 g507 (.n_ena(w249), .a(w256), .x(w257) );
	dmg_notif0 g508 (.n_ena(w249), .a(w700), .x(w259) );
	dmg_notif0 g509 (.n_ena(w249), .a(w853), .x(w310) );
	dmg_notif0 g510 (.n_ena(w249), .a(w250), .x(w66) );
	dmg_notif0 g511 (.n_ena(w170), .a(w319), .x(w318) );
	dmg_notif0 g512 (.n_ena(w62), .a(w458), .x(w567) );
	dmg_notif0 g513 (.n_ena(w140), .a(w527), .x(w460) );
	dmg_notif0 g514 (.n_ena(w140), .a(w901), .x(w168) );
	dmg_notif0 g515 (.n_ena(w140), .a(w901), .x(w59) );
	dmg_notif0 g516 (.n_ena(w140), .a(w527), .x(w60) );
	dmg_notif0 g517 (.n_ena(w140), .a(w526), .x(w63) );
	dmg_notif0 g518 (.n_ena(w140), .a(w526), .x(w9) );
	dmg_notif0 g519 (.n_ena(w140), .a(w534), .x(w141) );
	dmg_notif0 g520 (.n_ena(w140), .a(w534), .x(w178) );
	dmg_notif0 g521 (.n_ena(w140), .a(w558), .x(w465) );
	dmg_notif0 g522 (.n_ena(w140), .a(w558), .x(w567) );
	dmg_notif0 g523 (.n_ena(w140), .a(w561), .x(w164) );
	dmg_notif0 g524 (.n_ena(w140), .a(w561), .x(w5) );
	dmg_not g525 (.a(w603), .x(w64) );
	dmg_not g526 (.a(w47), .x(w129) );
	dmg_const g527 (.q0(w69), .q1(w149) );
	dmg_not2 g528 (.a(w560), .x(w392) );
	dmg_not2 g529 (.a(w138), .x(w137) );
	dmg_not2 g530 (.a(w138), .x(w62) );
	dmg_not2 g531 (.a(w889), .x(w123) );
	dmg_not2 g532 (.a(w3), .x(w518) );
	dmg_not2 g533 (.a(w912), .x(w170) );
	dmg_not2 g534 (.a(w697), .x(w37) );
	dmg_not2 g535 (.a(w391), .x(w390) );
	dmg_not2 g536 (.a(w399), .x(w427) );
	dmg_not2 g537 (.a(w860), .x(w569) );
	dmg_not2 g538 (.a(w188), .x(w189) );
	dmg_not2 g539 (.a(w713), .x(w409) );
	dmg_not2 g540 (.a(w104), .x(w79) );
	dmg_not2 g541 (.a(w230), .x(w229) );
	dmg_not2 g542 (.a(w96), .x(w95) );
	dmg_not2 g543 (.a(w423), .x(w424) );
	dmg_not2 g544 (.a(w200), .x(w44) );
	dmg_not2 g545 (.a(w57), .x(w58) );
	dmg_not2 g546 (.a(w210), .x(w209) );
	dmg_not2 g547 (.a(w492), .x(w491) );
	dmg_not2 g548 (.a(w162), .x(w11) );
	dmg_not2 g549 (.a(w551), .x(w140) );
	dmg_not2 g550 (.a(w765), .x(w576) );
	dmg_not2 g551 (.a(w617), .x(w304) );
	dmg_not2 g552 (.a(w634), .x(w249) );
	dmg_not2 g553 (.a(w378), .x(w635) );
	dmg_not2 g554 (.a(w820), .x(w245) );
	dmg_not2 g555 (.a(w842), .x(w179) );
	dmg_not2 g556 (.a(w557), .x(w556) );
	dmg_not2 g557 (.a(w126), .x(w127) );
	dmg_not2 g558 (.a(w564), .x(w563) );
	dmg_not2 g559 (.a(w491), .x(w648) );
	dmg_not2 g560 (.a(w509), .x(w177) );
	dmg_not2 g561 (.a(w114), .x(w113) );
	dmg_not2 g562 (.a(w336), .x(w290) );
	dmg_not2 g563 (.a(w370), .x(w280) );
	dmg_not2 g564 (.a(w339), .x(w274) );
	dmg_not2 g565 (.a(w23), .x(w330) );
	dmg_not2 g566 (.a(w758), .x(w28) );
	dmg_not2 g567 (.a(w852), .x(w223) );
	dmg_not2 g568 (.a(w455), .x(w403) );
	dmg_not2 g569 (.a(w160), .x(w637) );
	dmg_not2 g570 (.a(w406), .x(w183) );
	dmg_not g571 (.a(w225), .x(w226) );
	dmg_notif0 g572 (.n_ena(w170), .a(w910), .x(w52) );
	dmg_not g573 (.a(w98), .x(w99) );
	dmg_and g574 (.a(w454), .b(w888), .x(w206) );
	dmg_and g575 (.a(w4), .b(w101), .x(w102) );
	dmg_and g576 (.a(w101), .b(w100), .x(w3) );
	dmg_and g577 (.a(w2), .b(w205), .x(w532) );
	dmg_and g578 (.a(w2), .b(w1), .x(w204) );
	dmg_and g579 (.a(w1), .b(w393), .x(w144) );
	dmg_and g580 (.a(w208), .b(w4), .x(w53) );
	dmg_and g581 (.a(w53), .b(w54), .x(w332) );
	dmg_and g582 (.a(w857), .b(w155), .x(w154) );
	dmg_and g583 (.a(w858), .b(w857), .x(w406) );
	dmg_and g584 (.a(w408), .b(w407), .x(w792) );
	dmg_not g585 (.a(w863), .x(w508) );
	dmg_notif0 g586 (.n_ena(w635), .a(w849), .x(w279) );
	dmg_fa g587 (.cin(w813), .a(w104), .b(w103), .s(w533) );
	dmg_fa g588 (.cin(w810), .a(w188), .b(w187), .s(w448), .cout(w449) );
	dmg_fa g589 (.cin(w856), .a(w399), .b(w400), .cout(w699) );
	dmg_fa g590 (.cin(w181), .a(w105), .b(w519), .s(w182) );
	dmg_fa g591 (.cin(w523), .a(w447), .b(w522), .s(w180), .cout(w181) );
	dmg_fa g592 (.cin(w809), .a(w539), .b(w538), .s(w467), .cout(w466) );
	dmg_fa g593 (.cin(w151), .a(w398), .b(w805), .s(w150), .cout(w809) );
	dmg_fa g594 (.cin(w807), .a(w439), .b(w440), .s(w152), .cout(w151) );
	dmg_fa g595 (.cin(w69), .a(w388), .b(w387), .s(w68), .cout(w848) );
	dmg_fa g596 (.cin(w848), .a(w312), .b(w313), .s(w543), .cout(w542) );
	dmg_fa g597 (.cin(w541), .a(w540), .b(w110), .s(w479), .cout(w478) );
	dmg_fa g598 (.cin(w478), .a(w472), .b(w119), .s(w473), .cout(w477) );
	dmg_fa g599 (.cin(w711), .a(w446), .b(w445), .s(w485), .cout(w486) );
	dmg_fa g600 (.cin(w486), .a(w106), .b(w395), .s(w482), .cout(w481) );
	dmg_fa g601 (.cin(w477), .a(w316), .b(w315), .s(w476), .cout(w711) );
	dmg_fa g602 (.cin(w542), .a(w397), .b(w396), .s(w438), .cout(w541) );
	dmg_fa g603 (.cin(w466), .a(w471), .b(w470), .s(w468), .cout(w696) );
	dmg_fa g604 (.cin(w696), .a(w317), .b(w535), .s(w524), .cout(w523) );
	dmg_fa g605 (.cin(w903), .a(w200), .b(w201), .s(w812), .cout(w813) );
	dmg_fa g606 (.cin(w449), .a(w697), .b(w8), .s(w814), .cout(w903) );
	dmg_fa g607 (.cin(w699), .a(w230), .b(w231), .s(w698), .cout(w810) );
	dmg_fa g608 (.cin(w793), .a(w96), .b(w156), .cout(w856) );
	dmg_dffr g609 (.clk(w459), .nr1(w712), .d(w98), .nr2(w712), .q(w909) );
	dmg_dffr g610 (.clk(w833), .nr1(w410), .d(w714), .nr2(w410), .nq(w714), .q(w220) );
	dmg_dffr g611 (.clk(w199), .nr1(w371), .d(w758), .nr2(w371), .q(w373) );
	dmg_dffr g612 (.clk(w492), .nr1(w712), .d(w792), .nr2(w712), .q(w98) );
	dmg_dffr g613 (.clk(w492), .nr1(w712), .d(w100), .nr2(w712), .nq(w210) );
	dmg_dffr g614 (.clk(w495), .nr1(w650), .d(w881), .nr2(w650), .nq(w881), .q(w640) );
	dmg_dffr g615 (.clk(w199), .nr1(w371), .d(w23), .nr2(w371), .q(w338) );
	dmg_dffr g616 (.clk(w199), .nr1(w371), .d(w336), .nr2(w371), .q(w198) );
	dmg_dffr g617 (.clk(w199), .nr1(w371), .d(w339), .nr2(w371), .q(w331) );
	dmg_dffr g618 (.clk(w199), .nr1(w371), .d(w378), .nr2(w371), .q(w836) );
	dmg_dffr g619 (.clk(w707), .nr1(w650), .d(w495), .nr2(w650), .nq(w495), .q(w494) );
	dmg_dffr g620 (.clk(w199), .nr1(w371), .d(w634), .nr2(w371), .q(w693) );
	dmg_dffr g621 (.clk(w647), .nr1(w650), .d(w651), .nr2(w650), .nq(w651), .q(w517) );
	dmg_dffr g622 (.clk(w199), .nr1(w371), .d(w820), .nr2(w371), .q(w364) );
	dmg_dffr g623 (.clk(w199), .nr1(w371), .d(w765), .nr2(w371), .q(w379) );
	dmg_dffr g624 (.clk(w199), .nr1(w371), .d(w617), .nr2(w371), .q(w755) );
	dmg_dffr g625 (.clk(w651), .nr1(w650), .d(w707), .nr2(w650), .nq(w707), .q(w516) );
	dmg_dffr g626 (.clk(w710), .nr1(w650), .d(w806), .nr2(w650), .nq(w806), .q(w708) );
	dmg_dffr g627 (.clk(w881), .nr1(w650), .d(w710), .nr2(w650), .nq(w710), .q(w709) );
	dmg_dffr g628 (.clk(w199), .nr1(w371), .d(w370), .nr2(w371), .q(w756) );
	dmg_dffr g629 (.clk(w835), .nr1(w410), .d(w411), .nr2(w410), .nq(w411), .q(w219) );
	dmg_dffr g630 (.clk(w391), .nr1(w571), .d(w223), .nr2(w571), .q(w572) );
	dmg_dffr g631 (.clk(w390), .nr1(w252), .d(w791), .nr2(w252), .q(w254) );
	dmg_dffr g632 (.clk(w492), .nr1(w252), .d(w493), .nr2(w252), .nq(w855), .q(w791) );
	dmg_dffr g633 (.clk(w714), .nr1(w410), .d(w835), .nr2(w410), .nq(w835), .q(w574) );
	dmg_dffr g634 (.clk(w834), .nr1(w410), .d(w833), .nr2(w410), .nq(w833), .q(w575) );
	dmg_latchr_comp g635 (.n_ena(w227), .d(w594), .ena(w747), .nres(w372), .q(w897) );
	dmg_latchr_comp g636 (.n_ena(w227), .d(w413), .ena(w747), .nres(w372), .q(w789) );
	dmg_latchr_comp g637 (.n_ena(w295), .d(w433), .ena(w296), .nres(w787), .q(w796) );
	dmg_latchr_comp g638 (.n_ena(w295), .d(w594), .ena(w296), .nres(w787), .q(w861) );
	dmg_latchr_comp g639 (.n_ena(w443), .d(w402), .ena(w159), .nres(w11), .q(w400), .nq(w401) );
	dmg_latchr_comp g640 (.n_ena(w443), .d(w7), .ena(w159), .nres(w11), .q(w201), .nq(w202) );
	dmg_latchr_comp g641 (.n_ena(w443), .d(w6), .ena(w159), .nres(w11), .q(w8), .nq(w442) );
	dmg_latchr_comp g642 (.n_ena(w432), .d(w325), .ena(w437), .nres(w386), .q(w893) );
	dmg_latchr_comp g643 (.n_ena(w432), .d(w294), .ena(w437), .nres(w386), .q(w425) );
	dmg_latchr_comp g644 (.n_ena(w432), .d(w431), .ena(w437), .nres(w386), .q(w846) );
	dmg_latchr_comp g645 (.n_ena(w432), .d(w415), .ena(w437), .nres(w386), .q(w426) );
	dmg_latchr_comp g646 (.n_ena(w432), .d(w590), .ena(w437), .nres(w386), .q(w385) );
	dmg_latchr_comp g647 (.n_ena(w265), .d(w590), .ena(w90), .nres(w82), .q(w872) );
	dmg_latchr_comp g648 (.n_ena(w265), .d(w413), .ena(w90), .nres(w82), .q(w260) );
	dmg_latchr_comp g649 (.n_ena(w265), .d(w433), .ena(w90), .nres(w82), .q(w764) );
	dmg_latchr_comp g650 (.n_ena(w293), .d(w590), .ena(w40), .nres(w39), .q(w41) );
	dmg_latchr_comp g651 (.n_ena(w293), .d(w433), .ena(w40), .nres(w39), .q(w38) );
	dmg_latchr_comp g652 (.n_ena(w293), .d(w431), .ena(w40), .nres(w39), .q(w430) );
	dmg_latchr_comp g653 (.n_ena(w265), .d(w294), .ena(w90), .nres(w82), .q(w83) );
	dmg_latchr_comp g654 (.n_ena(w265), .d(w325), .ena(w90), .nres(w82), .q(w91) );
	dmg_latchr_comp g655 (.n_ena(w265), .d(w415), .ena(w90), .nres(w82), .q(w94) );
	dmg_latchr_comp g656 (.n_ena(w265), .d(w431), .ena(w90), .nres(w82), .q(w89) );
	dmg_latchr_comp g657 (.n_ena(w184), .d(w234), .ena(w10), .nres(w11), .q(w639), .nq(w638) );
	dmg_latchr_comp g658 (.n_ena(w443), .d(w12), .ena(w159), .nres(w11), .q(w231), .nq(w232) );
	dmg_latchr_comp g659 (.n_ena(w350), .d(w415), .ena(w414), .nres(w351), .q(w357) );
	dmg_latchr_comp g660 (.n_ena(w350), .d(w325), .ena(w414), .nres(w351), .q(w782) );
	dmg_latchr_comp g661 (.n_ena(w350), .d(w294), .ena(w414), .nres(w351), .q(w882) );
	dmg_latchr_comp g662 (.n_ena(w350), .d(w431), .ena(w414), .nres(w351), .q(w781) );
	dmg_latchr_comp g663 (.n_ena(w350), .d(w413), .ena(w414), .nres(w351), .q(w907) );
	dmg_latchr_comp g664 (.n_ena(w583), .d(w325), .ena(w585), .nres(w584), .q(w627) );
	dmg_latchr_comp g665 (.n_ena(w583), .d(w415), .ena(w585), .nres(w584), .q(w602) );
	dmg_latchr_comp g666 (.d(w294), .ena(w585), .nres(w584), .q(w744), .n_ena(w583) );
	dmg_latchr_comp g667 (.n_ena(w583), .d(w431), .ena(w585), .nres(w584), .q(w689) );
	dmg_latchr_comp g668 (.n_ena(w591), .d(w431), .ena(w77), .nres(w593), .q(w676) );
	dmg_latchr_comp g669 (.n_ena(w591), .d(w594), .ena(w77), .nres(w593), .q(w78) );
	dmg_latchr_comp g670 (.n_ena(w369), .d(w594), .ena(w512), .nres(w21), .q(w612) );
	dmg_latchr_comp g671 (.n_ena(w369), .d(w433), .ena(w512), .nres(w21), .q(w588) );
	dmg_latchr_comp g672 (.n_ena(w369), .d(w294), .ena(w512), .nres(w21), .q(w771) );
	dmg_latchr_comp g673 (.n_ena(w369), .d(w415), .ena(w512), .nres(w21), .q(w20) );
	dmg_latchr_comp g674 (.n_ena(w369), .d(w431), .ena(w512), .nres(w21), .q(w608) );
	dmg_latchr_comp g675 (.n_ena(w591), .d(w433), .ena(w77), .nres(w593), .q(w587) );
	dmg_latchr_comp g676 (.n_ena(w591), .d(w415), .ena(w77), .nres(w593), .q(w604) );
	dmg_latchr_comp g677 (.n_ena(w595), .d(w433), .ena(w600), .nres(w362), .q(w672) );
	dmg_latchr_comp g678 (.n_ena(w595), .d(w413), .ena(w600), .nres(w362), .q(w845) );
	dmg_latchr_comp g679 (.n_ena(w595), .d(w590), .ena(w600), .nres(w362), .q(w626) );
	dmg_latchr_comp g680 (.n_ena(w595), .d(w594), .ena(w600), .nres(w362), .q(w361) );
	dmg_latchr_comp g681 (.n_ena(w583), .d(w433), .ena(w585), .nres(w584), .q(w586) );
	dmg_latchr_comp g682 (.n_ena(w583), .d(w590), .ena(w585), .nres(w584), .q(w629) );
	dmg_latchr_comp g683 (.n_ena(w583), .d(w413), .ena(w585), .nres(w584), .q(w628) );
	dmg_latchr_comp g684 (.n_ena(w583), .d(w594), .ena(w585), .nres(w584), .q(w740) );
	dmg_latchr_comp g685 (.n_ena(w595), .d(w431), .ena(w600), .nres(w362), .q(w774) );
	dmg_latchr_comp g686 (.n_ena(w595), .d(w325), .ena(w600), .nres(w362), .q(w599) );
	dmg_latchr_comp g687 (.n_ena(w595), .d(w294), .ena(w600), .nres(w362), .q(w596) );
	dmg_latchr_comp g688 (.n_ena(w595), .d(w415), .ena(w600), .nres(w362), .q(w601) );
	dmg_latchr_comp g689 (.n_ena(w591), .d(w325), .ena(w77), .nres(w593), .q(w605) );
	dmg_latchr_comp g690 (.n_ena(w591), .d(w413), .ena(w77), .nres(w593), .q(w76) );
	dmg_latchr_comp g691 (.n_ena(w369), .d(w325), .ena(w512), .nres(w21), .q(w611) );
	dmg_latchr_comp g692 (.n_ena(w369), .d(w413), .ena(w512), .nres(w21), .q(w368) );
	dmg_latchr_comp g693 (.n_ena(w369), .d(w590), .ena(w512), .nres(w21), .q(w592) );
	dmg_latchr_comp g694 (.n_ena(w591), .d(w590), .ena(w77), .nres(w593), .q(w71) );
	dmg_latchr_comp g695 (.n_ena(w591), .d(w294), .ena(w77), .nres(w593), .q(w678) );
	dmg_latchr_comp g696 (.n_ena(w350), .d(w433), .ena(w414), .nres(w351), .q(w353) );
	dmg_latchr_comp g697 (.n_ena(w350), .d(w594), .ena(w414), .nres(w351), .q(w352) );
	dmg_latchr_comp g698 (.n_ena(w350), .d(w590), .ena(w414), .nres(w351), .q(w356) );
	dmg_latchr_comp g699 (.n_ena(w184), .d(w7), .ena(w10), .nres(w11), .q(w522), .nq(w528) );
	dmg_latchr_comp g700 (.n_ena(w184), .d(w521), .ena(w10), .nres(w11), .q(w519), .nq(w520) );
	dmg_latchr_comp g701 (.n_ena(w184), .d(w12), .ena(w10), .nres(w11), .q(w538), .nq(w537) );
	dmg_latchr_comp g702 (.n_ena(w184), .d(w6), .ena(w10), .nres(w11), .q(w535), .nq(w536) );
	dmg_latchr_comp g703 (.n_ena(w184), .d(w402), .ena(w10), .nres(w11), .q(w805), .nq(w441) );
	dmg_latchr_comp g704 (.n_ena(w184), .d(w158), .ena(w10), .nres(w11), .q(w440), .nq(w646) );
	dmg_latchr_comp g705 (.n_ena(w432), .d(w413), .ena(w437), .nres(w386), .q(w799) );
	dmg_latchr_comp g706 (.n_ena(w432), .d(w594), .ena(w437), .nres(w386), .q(w800) );
	dmg_latchr_comp g707 (.n_ena(w432), .d(w433), .ena(w437), .nres(w386), .q(w801) );
	dmg_latchr_comp g708 (.n_ena(w227), .d(w325), .ena(w747), .nres(w372), .q(w783) );
	dmg_latchr_comp g709 (.n_ena(w227), .d(w415), .ena(w747), .nres(w372), .q(w374) );
	dmg_latchr_comp g710 (.n_ena(w227), .d(w294), .ena(w747), .nres(w372), .q(w751) );
	dmg_latchr_comp g711 (.n_ena(w227), .d(w431), .ena(w747), .nres(w372), .q(w380) );
	dmg_latchr_comp g712 (.n_ena(w265), .d(w594), .ena(w90), .nres(w82), .q(w264) );
	dmg_latchr_comp g713 (.n_ena(w293), .d(w325), .ena(w40), .nres(w39), .q(w416) );
	dmg_latchr_comp g714 (.n_ena(w293), .d(w415), .ena(w40), .nres(w39), .q(w434) );
	dmg_latchr_comp g715 (.n_ena(w293), .d(w294), .ena(w40), .nres(w39), .q(w615) );
	dmg_latchr_comp g716 (.n_ena(w293), .d(w413), .ena(w40), .nres(w39), .q(w412) );
	dmg_latchr_comp g717 (.n_ena(w293), .d(w594), .ena(w40), .nres(w39), .q(w196) );
	dmg_latchr_comp g718 (.n_ena(w227), .d(w433), .ena(w747), .nres(w372), .q(w730) );
	dmg_latchr_comp g719 (.n_ena(w295), .d(w294), .ena(w296), .nres(w787), .q(w759) );
	dmg_latchr_comp g720 (.n_ena(w295), .d(w325), .ena(w296), .nres(w787), .q(w760) );
	dmg_latchr_comp g721 (.n_ena(w295), .d(w415), .ena(w296), .nres(w787), .q(w762) );
	dmg_latchr_comp g722 (.n_ena(w227), .d(w590), .ena(w747), .nres(w372), .q(w790) );
	dmg_latchr_comp g723 (.n_ena(w295), .d(w431), .ena(w296), .nres(w787), .q(w228) );
	dmg_latchr_comp g724 (.n_ena(w295), .d(w590), .ena(w296), .nres(w787), .q(w36) );
	dmg_latchr_comp g725 (.n_ena(w295), .d(w413), .ena(w296), .nres(w787), .q(w788) );
	dmg_latchr_comp g726 (.n_ena(w184), .d(w185), .ena(w10), .nres(w11), .q(w470), .nq(w469) );
	dmg_latchr_comp g727 (.n_ena(w443), .d(w234), .ena(w159), .nres(w11), .q(w422), .nq(w864) );
	dmg_latchr_comp g728 (.n_ena(w443), .d(w158), .ena(w159), .nres(w11), .q(w156), .nq(w157) );
	dmg_latchr_comp g729 (.n_ena(w443), .d(w185), .ena(w159), .nres(w11), .q(w187), .nq(w186) );
	dmg_latchr_comp g730 (.n_ena(w443), .d(w521), .ena(w159), .nres(w11), .q(w103), .nq(w890) );
	dmg_notif0 g731 (.n_ena(w170), .a(w396), .x(w133) );
	dmg_not g732 (.a(w218), .x(w269) );
	dmg_latch g733 (.ena(w165), .d(w164), .q(w175), .nq(w176) );
	dmg_latch g734 (.ena(w165), .d(w59), .q(w905), .nq(w496) );
	dmg_latch g735 (.ena(w165), .d(w5), .q(w241), .nq(w238) );
	dmg_latch g736 (.ena(w165), .d(w510), .q(w505), .nq(w504) );
	dmg_latch g737 (.ena(w165), .d(w168), .q(w705), .nq(w704) );
	dmg_latch g738 (.ena(w165), .d(w465), .q(w14), .nq(w13) );
	dmg_latch g739 (.ena(w165), .d(w63), .q(w121), .nq(w122) );
	dmg_latch g740 (.ena(w165), .d(w178), .q(w566), .nq(w565) );
	dmg_latch g741 (.ena(w165), .d(w60), .q(w501), .nq(w706) );
	dmg_latch g742 (.ena(w165), .d(w460), .q(w461), .nq(w462) );
	dmg_latch g743 (.ena(w165), .d(w169), .q(w236), .nq(w235) );
	dmg_latch g744 (.ena(w165), .d(w9), .q(w502), .nq(w503) );
	dmg_latch g745 (.ena(w165), .d(w567), .q(w240), .nq(w239) );
	dmg_latch g746 (.ena(w165), .d(w163), .q(w506), .nq(w507) );
	dmg_latch g747 (.ena(w165), .d(w243), .q(w111), .nq(w112) );
	dmg_latch g748 (.ena(w165), .d(w141), .q(w420), .nq(w421) );
	dmg_bufif0 g749 (.a0(w112), .n_ena(w113), .a1(w112), .x(w12) );
	dmg_bufif0 g750 (.a0(w239), .n_ena(w113), .a1(w239), .x(w7) );
	dmg_bufif0 g751 (.a0(w462), .n_ena(w113), .a1(w462), .x(w158) );
	dmg_bufif0 g752 (.a0(w507), .n_ena(w177), .a1(w507), .x(w12) );
	dmg_bufif0 g753 (.a0(w421), .n_ena(w177), .a1(w421), .x(w185) );
	dmg_bufif0 g754 (.a0(w503), .n_ena(w177), .a1(w503), .x(w402) );
	dmg_bufif0 g755 (.a0(w504), .n_ena(w177), .a1(w504), .x(w234) );
	dmg_bufif0 g756 (.a0(w706), .n_ena(w177), .a1(w706), .x(w158) );
	dmg_bufif0 g757 (.a0(w13), .n_ena(w177), .a1(w13), .x(w7) );
	dmg_bufif0 g758 (.a0(w565), .n_ena(w113), .a1(w565), .x(w185) );
	dmg_bufif0 g759 (.a0(w704), .n_ena(w113), .a1(w704), .x(w521) );
	dmg_bufif0 g760 (.a0(w238), .n_ena(w113), .a1(w238), .x(w6) );
	dmg_bufif0 g761 (.a0(w122), .n_ena(w113), .a1(w122), .x(w402) );
	dmg_bufif0 g762 (.a0(w235), .n_ena(w113), .a1(w235), .x(w234) );
	dmg_bufif0 g763 (.a0(w496), .n_ena(w177), .a1(w496), .x(w521) );
	dmg_bufif0 g764 (.a0(w176), .n_ena(w177), .a1(w176), .x(w6) );
	dmg_xor g765 (.a(w258), .b(w66), .x(w319) );
	dmg_xor g766 (.a(w36), .b(w44), .x(w35) );
	dmg_xor g767 (.a(w790), .b(w44), .x(w854) );
	dmg_xor g768 (.a(w788), .b(w189), .x(w795) );
	dmg_xor g769 (.a(w730), .b(w37), .x(w731) );
	dmg_xor g770 (.a(w196), .b(w79), .x(w195) );
	dmg_xor g771 (.a(w412), .b(w189), .x(w679) );
	dmg_xor g772 (.a(w760), .b(w95), .x(w30) );
	dmg_xor g773 (.a(w759), .b(w424), .x(w31) );
	dmg_xor g774 (.a(w762), .b(w427), .x(w29) );
	dmg_xor g775 (.a(w228), .b(w229), .x(w749) );
	dmg_xor g776 (.a(w801), .b(w37), .x(w797) );
	dmg_xor g777 (.a(w800), .b(w79), .x(w383) );
	dmg_xor g778 (.a(w799), .b(w189), .x(w798) );
	dmg_xor g779 (.a(w783), .b(w95), .x(w784) );
	dmg_xor g780 (.a(w374), .b(w427), .x(w375) );
	dmg_xor g781 (.a(w380), .b(w229), .x(w376) );
	dmg_xor g782 (.a(w751), .b(w424), .x(w785) );
	dmg_xor g783 (.a(w83), .b(w424), .x(w84) );
	dmg_xor g784 (.a(w89), .b(w229), .x(w88) );
	dmg_xor g785 (.a(w94), .b(w427), .x(w93) );
	dmg_xor g786 (.a(w91), .b(w95), .x(w92) );
	dmg_xor g787 (.a(w71), .b(w44), .x(w72) );
	dmg_xor g788 (.a(w678), .b(w424), .x(w677) );
	dmg_xor g789 (.a(w596), .b(w424), .x(w597) );
	dmg_xor g790 (.a(w601), .b(w427), .x(w745) );
	dmg_xor g791 (.a(w356), .b(w44), .x(w355) );
	dmg_xor g792 (.a(w353), .b(w37), .x(w354) );
	dmg_xor g793 (.a(w352), .b(w79), .x(w780) );
	dmg_xor g794 (.a(w586), .b(w37), .x(w191) );
	dmg_xor g795 (.a(w740), .b(w79), .x(w742) );
	dmg_xor g796 (.a(w629), .b(w44), .x(w741) );
	dmg_xor g797 (.a(w628), .b(w189), .x(w192) );
	dmg_xor g798 (.a(w626), .b(w44), .x(w625) );
	dmg_xor g799 (.a(w672), .b(w37), .x(w884) );
	dmg_xor g800 (.a(w845), .b(w189), .x(w883) );
	dmg_xor g801 (.a(w361), .b(w79), .x(w360) );
	dmg_xor g802 (.a(w605), .b(w95), .x(w606) );
	dmg_xor g803 (.a(w599), .b(w95), .x(w598) );
	dmg_xor g804 (.a(w774), .b(w229), .x(w773) );
	dmg_xor g805 (.a(w604), .b(w427), .x(w607) );
	dmg_xor g806 (.a(w76), .b(w189), .x(w75) );
	dmg_xor g807 (.a(w587), .b(w37), .x(w74) );
	dmg_xor g808 (.a(w78), .b(w79), .x(w73) );
	dmg_xor g809 (.a(w611), .b(w95), .x(w610) );
	dmg_xor g810 (.a(w608), .b(w229), .x(w18) );
	dmg_xor g811 (.a(w20), .b(w427), .x(w19) );
	dmg_xor g812 (.a(w771), .b(w424), .x(w609) );
	dmg_xor g813 (.a(w612), .b(w79), .x(w80) );
	dmg_xor g814 (.a(w588), .b(w37), .x(w366) );
	dmg_xor g815 (.a(w676), .b(w229), .x(w673) );
	dmg_xor g816 (.a(w907), .b(w189), .x(w908) );
	dmg_xor g817 (.a(w781), .b(w229), .x(w777) );
	dmg_xor g818 (.a(w782), .b(w95), .x(w359) );
	dmg_xor g819 (.a(w357), .b(w427), .x(w358) );
	dmg_xor g820 (.a(w882), .b(w424), .x(w671) );
	dmg_xor g821 (.a(w602), .b(w427), .x(w190) );
	dmg_xor g822 (.a(w744), .b(w424), .x(w670) );
	dmg_xor g823 (.a(w689), .b(w229), .x(w614) );
	dmg_xor g824 (.a(w627), .b(w95), .x(w669) );
	dmg_xor g825 (.a(w258), .b(w257), .x(w754) );
	dmg_xor g826 (.a(w592), .b(w44), .x(w81) );
	dmg_xor g827 (.a(w368), .b(w189), .x(w367) );
	dmg_xor g828 (.a(w434), .b(w427), .x(w428) );
	dmg_xor g829 (.a(w615), .b(w424), .x(w418) );
	dmg_xor g830 (.a(w430), .b(w229), .x(w429) );
	dmg_xor g831 (.a(w416), .b(w95), .x(w417) );
	dmg_xor g832 (.a(w893), .b(w95), .x(w255) );
	dmg_xor g833 (.a(w425), .b(w424), .x(w435) );
	dmg_xor g834 (.a(w846), .b(w229), .x(w436) );
	dmg_xor g835 (.a(w426), .b(w427), .x(w847) );
	dmg_xor g836 (.a(w385), .b(w44), .x(w384) );
	dmg_xor g837 (.a(w260), .b(w189), .x(w261) );
	dmg_xor g838 (.a(w764), .b(w37), .x(w262) );
	dmg_xor g839 (.a(w872), .b(w44), .x(w763) );
	dmg_xor g840 (.a(w38), .b(w37), .x(w43) );
	dmg_xor g841 (.a(w41), .b(w44), .x(w42) );
	dmg_xor g842 (.a(w897), .b(w79), .x(w898) );
	dmg_xor g843 (.a(w789), .b(w189), .x(w732) );
	dmg_xor g844 (.a(w861), .b(w79), .x(w34) );
	dmg_xor g845 (.a(w796), .b(w37), .x(w794) );
	dmg_xor g846 (.a(w258), .b(w259), .x(w910) );
	dmg_xor g847 (.a(w258), .b(w310), .x(w911) );
	dmg_or g848 (.a(w223), .b(w224), .x(w225) );
	dmg_or g849 (.a(w223), .b(w346), .x(w345) );
	dmg_or g850 (.a(w223), .b(w217), .x(w216) );
	dmg_or g851 (.a(w223), .b(w268), .x(w267) );
	dmg_or g852 (.a(w223), .b(w271), .x(w322) );
	dmg_or g853 (.a(w573), .b(w572), .x(w834) );
	dmg_or g854 (.a(w27), .b(w373), .x(w894) );
	dmg_or g855 (.a(w223), .b(w222), .x(w616) );
	dmg_or g856 (.a(w223), .b(w665), .x(w913) );
	dmg_or g857 (.a(w27), .b(w338), .x(w70) );
	dmg_or g858 (.a(w822), .b(w69), .x(w752) );
	dmg_or g859 (.a(w334), .b(w335), .x(w377) );
	dmg_or g860 (.a(w803), .b(w24), .x(w25) );
	dmg_or g861 (.a(w27), .b(w836), .x(w837) );
	dmg_or g862 (.a(w27), .b(w755), .x(w26) );
	dmg_or g863 (.a(w630), .b(w25) );
	dmg_or g864 (.a(w109), .b(w479), .x(w480) );
	dmg_or g865 (.a(w493), .b(w492), .x(w647) );
	dmg_or g866 (.a(w821), .b(w621), .x(w620) );
	dmg_or g867 (.a(w223), .b(w660), .x(w661) );
	dmg_or g868 (.a(w223), .b(w514), .x(w513) );
	dmg_or g869 (.a(w27), .b(w364), .x(w363) );
	dmg_or g870 (.a(w27), .b(w693), .x(w692) );
	dmg_or g871 (.a(w622), .b(w619), .x(w618) );
	dmg_or g872 (.a(w786), .b(w377), .x(w621) );
	dmg_or g873 (.a(w766), .b(w620), .x(w619) );
	dmg_or g874 (.a(w802), .b(w618), .x(w24) );
	dmg_or g875 (.a(w804), .b(w767), .x(w545) );
	dmg_or g876 (.a(w753), .b(w752), .x(w335) );
	dmg_or g877 (.a(w27), .b(w379), .x(w337) );
	dmg_or g878 (.a(w27), .b(w198), .x(w197) );
	dmg_or g879 (.a(w27), .b(w331), .x(w22) );
	dmg_or g880 (.a(w27), .b(w756), .x(w757) );
	dmg_or g881 (.a(w223), .b(w299), .x(w298) );
	dmg_or g882 (.a(w409), .b(w688), .x(w687) );
	dmg_or g883 (.a(w570), .b(w569), .x(w568) );
	dmg_and g884 (.a(w205), .b(w393), .x(w811) );
	dmg_and g885 (.a(w210), .b(w4), .x(w211) );
	dmg_and g886 (.a(w220), .b(w219), .x(w573) );
	dmg_and g887 (.a(w125), .b(w508), .x(w557) );
	dmg_and g888 (.a(w463), .b(w125), .x(w126) );
	dmg_nand4 g889 (.a(w300), .b(w301), .c(w221), .d(w218), .x(w514) );
	dmg_nand4 g890 (.a(w515), .b(w301), .c(w272), .d(w218), .x(w665) );
	dmg_nand4 g891 (.a(w515), .b(w301), .c(w221), .d(w218), .x(w222) );
	dmg_nand4 g892 (.a(w300), .b(w301), .c(w272), .d(w218), .x(w660) );
	dmg_nand4 g893 (.a(w515), .b(w270), .c(w221), .d(w269), .x(w346) );
	dmg_nand4 g894 (.a(w300), .b(w270), .c(w221), .d(w218), .x(w217) );
	dmg_nand4 g895 (.a(w300), .b(w270), .c(w221), .d(w269), .x(w268) );
	dmg_nand4 g896 (.a(w515), .b(w270), .c(w272), .d(w218), .x(w224) );
	dmg_nand4 g897 (.a(w515), .b(w270), .c(w221), .d(w218), .x(w299) );
	dmg_nand4 g898 (.a(w300), .b(w270), .c(w272), .d(w218), .x(w271) );
	dmg_nor4 g899 (.a(w679), .b(w43), .c(w42), .d(w195), .x(w194) );
	dmg_nor4 g900 (.a(w418), .b(w417), .c(w428), .d(w429), .x(w193) );
	dmg_nor4 g901 (.a(w261), .b(w262), .c(w763), .d(w263), .x(w86) );
	dmg_xor g902 (.a(w264), .b(w79), .x(w263) );
	dmg_nor4 g903 (.a(w84), .b(w92), .c(w93), .d(w88), .x(w87) );
	dmg_nor4 g904 (.a(w367), .b(w366), .c(w81), .d(w80), .x(w16) );
	dmg_nor4 g905 (.a(w609), .b(w610), .c(w19), .d(w18), .x(w17) );
	dmg_nor4 g906 (.a(w75), .b(w74), .c(w72), .d(w73), .x(w675) );
	dmg_nor4 g907 (.a(w597), .b(w598), .c(w745), .d(w773), .x(w775) );
	dmg_nor4 g908 (.a(w677), .b(w606), .c(w607), .d(w673), .x(w674) );
	dmg_nor4 g909 (.a(w908), .b(w354), .c(w355), .d(w780), .x(w779) );
	dmg_nor4 g910 (.a(w883), .b(w884), .c(w625), .d(w360), .x(w624) );
	dmg_nor4 g911 (.a(w671), .b(w359), .c(w358), .d(w777), .x(w778) );
	dmg_nor4 g912 (.a(w192), .b(w191), .c(w741), .d(w742), .x(w743) );
	dmg_nor4 g913 (.a(w670), .b(w669), .c(w190), .d(w614), .x(w613) );
	dmg_nor4 g914 (.a(w785), .b(w784), .c(w375), .d(w376), .x(w748) );
	dmg_nor4 g915 (.a(w31), .b(w30), .c(w29), .d(w749), .x(w32) );
	dmg_nor4 g916 (.a(w435), .b(w255), .c(w847), .d(w436), .x(w45) );
	dmg_nor4 g917 (.a(w795), .b(w794), .c(w35), .d(w34), .x(w33) );
	dmg_nor4 g918 (.a(w798), .b(w797), .c(w384), .d(w383), .x(w382) );
	dmg_nor4 g919 (.a(w732), .b(w731), .c(w854), .d(w898), .x(w761) );
	dmg_nand3 g920 (.a(w332), .b(w87), .c(w86), .x(w768) );
	dmg_nand3 g921 (.a(w332), .b(w193), .c(w194), .x(w333) );
	dmg_nand3 g922 (.a(w332), .b(w32), .c(w33), .x(w633) );
	dmg_nand3 g923 (.a(w332), .b(w748), .c(w761), .x(w750) );
	dmg_nand3 g924 (.a(w332), .b(w45), .c(w382), .x(w381) );
	dmg_nand3 g925 (.a(w332), .b(w613), .c(w743), .x(w631) );
	dmg_nand3 g926 (.a(w332), .b(w674), .c(w675), .x(w746) );
	dmg_nand3 g927 (.a(w332), .b(w17), .c(w16), .x(w365) );
	dmg_not g928 (.a(w419), .x(w413) );
	dmg_or3 g929 (.a(w254), .b(w253), .c(w855), .x(w860) );
	dmg_nor g930 (.a(w409), .b(w570), .x(w650) );
	dmg_nor g931 (.a(w333), .b(w335), .x(w336) );
	dmg_nor g932 (.a(w633), .b(w752), .x(w758) );
	dmg_nor g933 (.a(w768), .b(w24), .x(w23) );
	dmg_nor g934 (.a(w746), .b(w621), .x(w634) );
	dmg_nor g935 (.a(w365), .b(w69), .x(w339) );
	dmg_nor g936 (.a(w623), .b(w619), .x(w820) );
	dmg_not4 g937 (.a(w563), .x(w391) );
	dmg_dffrnq_comp g938 (.nr1(w149), .d(w130), .ck(w648), .cck(w491), .nr2(w149), .nq(w212) );
	dmg_dffrnq_comp g939 (.nr1(w149), .d(w555), .ck(w648), .cck(w491), .nr2(w149), .nq(w531) );
	dmg_dffrnq_comp g940 (.nr1(w149), .d(w128), .ck(w648), .cck(w491), .nr2(w149), .nq(w652) );
	dmg_dffrnq_comp g941 (.nr1(w149), .d(w129), .ck(w648), .cck(w491), .nr2(w149), .nq(w490) );
	dmg_dffrnq_comp g942 (.nr1(w149), .d(w147), .ck(w648), .cck(w491), .nr2(w149), .nq(w840) );
	dmg_dffrnq_comp g943 (.nr1(w149), .d(w148), .ck(w648), .cck(w491), .nr2(w149), .nq(w649) );
	dmg_and3 g944 (.a(w463), .b(w206), .c(w115), .x(w114) );
	dmg_and3 g945 (.a(w115), .b(w206), .c(w508), .x(w509) );
	dmg_aon g946 (.a0(w206), .a1(w205), .b(w124), .x(w125) );
	dmg_not4 g947 (.a(w392), .x(w1) );
	dmg_nand3 g948 (.a(w453), .b(w454), .c(w1), .x(w902) );
	dmg_aon22 g949 (.a0(w207), .a1(w206), .b0(w888), .b1(w456), .x(w889) );
	dmg_nor3 g950 (.a(w455), .b(w3), .c(w102), .x(w888) );
	dmg_or3 g951 (.a(w3), .b(w4), .c(w455), .x(w48) );
	dmg_oai g952 (.a0(w454), .a1(w455), .b(w548), .x(w547) );
	dmg_not4 g953 (.a(w637), .x(w205) );
	dmg_nor_latch g954 (.s(w98), .r(w568), .q(w100) );
	dmg_oan g955 (.a0(w909), .a1(w99), .b(w712), .x(w713) );
	dmg_nand3 g956 (.a(w547), .b(w546), .c(w56), .x(w57) );
	dmg_and3 g957 (.a(w815), .b(w209), .c(w816), .x(w852) );
	dmg_and3 g958 (.a(w167), .b(w172), .c(w902), .x(w166) );
	dmg_nand g959 (.a(w3), .b(w815), .x(w167) );
	dmg_nand g960 (.a(w3), .b(w55), .x(w56) );
	dmg_nand5 g961 (.a(w746), .b(w632), .c(w333), .d(w633), .e(w365), .x(w804) );
	dmg_nand5 g962 (.a(w631), .b(w768), .c(w381), .d(w623), .e(w750), .x(w767) );
	dmg_nor g963 (.a(w632), .b(w377), .x(w378) );
	dmg_nor g964 (.a(w631), .b(w25), .x(w370) );
	dmg_nor g965 (.a(w381), .b(w618), .x(w617) );
	dmg_aon22 g966 (.a0(w387), .a1(w818), .b0(w109), .b1(w754), .x(w695) );
	dmg_nand6 g967 (.a(w474), .b(w475), .c(w484), .d(w483), .e(w481), .f(w480), .x(w817) );
	dmg_nor g968 (.a(w750), .b(w620), .x(w765) );
	dmg_nand3 g969 (.a(w332), .b(w775), .c(w624), .x(w623) );
	dmg_nand3 g970 (.a(w332), .b(w778), .c(w779), .x(w632) );
	dmg_ha g971 (.a(w389), .b(w639), .cout(w807), .s(w808) );
	dmg_and4 g972 (.a(w517), .b(w516), .c(w708), .d(w494), .x(w493) );
	dmg_ha g973 (.a(w423), .b(w422), .cout(w793) );
endmodule // PPU2