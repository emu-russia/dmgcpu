// SM83 Decoder1.

module Decoder1 (a, d, clk);

	input wire [25:0] a;
	output wire [106:0] d;
	input wire clk;

endmodule // Decoder1
