
module Decoder1 (CLK2, a, d);

	input CLK2;
	input [25:0] a;
	output [106:0] d;

endmodule // Decoder1
