
module DataBridge( DataOut, DV, DL );

	input DataOut;
	input [7:0] DV;
	inout [7:0] DL;

endmodule // DataBridge
