module MMIO (  reset, clk2, clk4, osc_stable, clk_ena, osc_ena, clk6, clk9, n_reset2, cpu_wr_sync, cpu_m1, n_cpu_m1, 
	a, d, 
	cpu_irq_trig, cpu_irq_ack, cpu_rd, cpu_wr, 
	n_DRV_HIGH_a, n_INPUT_a, DRV_LOW_a, 
	n_DRV_HIGH_nrd, n_INPUT_nrd, DRV_LOW_nrd, n_DRV_HIGH_nwr, n_INPUT_nwr, DRV_LOW_nwr, n_t1_frompad, n_t2_frompad, CONST0, n_ena_pu_db, n_dma_phi, 
	dma_a, dma_a_15, dma_run, soc_wr, soc_rd, lfo_512Hz, ppu_rd, ppu_wr, int_serial, sc_read, sb_read, sc_write, n_sb_write, lfo_16384Hz, ppu_clk, vram_to_oam, non_vram_mreq, 
	test_1, test_2, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, n_test_reset, n_ext_addr_en, addr_latch, int_jp, FF60_D1, ffxx, n_ppu_hard_reset, ff46, dma_addr_ext, cpu_vram_oam_rd, oam_dma_wr, ppu_int_stat, ppu_int_vbl, clk6_delay);

	input wire reset;
	input wire clk2;
	input wire clk4;
	output wire osc_stable;
	input wire clk_ena;
	input wire osc_ena;
	input wire clk6;
	input wire clk9;
	input wire n_reset2;
	input wire cpu_wr_sync;
	input wire cpu_m1;
	output wire n_cpu_m1;
	inout wire [14:0] a; 			// a[15] is not used    ⚠️ bidir
	inout wire [7:0] d;
	output wire [4:0] cpu_irq_trig;
	input wire [4:0] cpu_irq_ack;
	input wire cpu_rd;
	input wire cpu_wr;
	output wire [14:8] n_DRV_HIGH_a;
	input wire [14:8] n_INPUT_a;
	output wire [14:8] DRV_LOW_a;
	output wire n_DRV_HIGH_nrd;
	input wire n_INPUT_nrd;
	output wire DRV_LOW_nrd;
	output wire n_DRV_HIGH_nwr;
	input wire n_INPUT_nwr;
	output wire DRV_LOW_nwr;
	input wire n_t1_frompad;
	input wire n_t2_frompad;
	inout wire CONST0;
	output wire n_ena_pu_db;
	output wire n_dma_phi;
	output wire [12:0] dma_a;
	output wire dma_a_15;
	output wire dma_run;
	output wire soc_wr;
	output wire soc_rd;
	output wire lfo_512Hz;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire int_serial;
	output wire sc_read;
	output wire sb_read;
	output wire sc_write;
	output wire n_sb_write;
	output wire lfo_16384Hz;
	input wire ppu_clk;
	output wire vram_to_oam;
	input wire non_vram_mreq;
	output wire test_1;
	output wire test_2;
	output wire n_extdb_to_intdb;
	output wire n_dblatch_to_intdb;
	output wire n_intdb_to_extdb;
	output wire n_test_reset;
	output wire n_ext_addr_en;
	output wire addr_latch;
	input wire int_jp;
	input wire FF60_D1;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ff46;
	output wire dma_addr_ext;
	output wire cpu_vram_oam_rd;
	output wire oam_dma_wr;
	input wire ppu_int_stat;
	input wire ppu_int_vbl;
	input wire clk6_delay;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;

	assign DRV_LOW_a[13] = w1;
	assign n_DRV_HIGH_a[13] = w7;
	assign w6 = n_INPUT_a[13];
	assign n_DRV_HIGH_a[12] = w51;
	assign DRV_LOW_a[12] = w289;
	assign n_DRV_HIGH_a[11] = w288;
	assign w233 = n_INPUT_a[8];
	assign n_DRV_HIGH_a[9] = w234;
	assign DRV_LOW_a[9] = w268;
	assign n_DRV_HIGH_a[8] = w291;
	assign DRV_LOW_a[8] = w292;
	assign w10 = n_INPUT_a[11];
	assign DRV_LOW_a[11] = w290;
	assign w267 = n_INPUT_a[9];
	assign w262 = clk_ena;
	assign w263 = n_INPUT_a[14];
	assign n_DRV_HIGH_a[14] = w265;
	assign DRV_LOW_a[14] = w266;
	assign osc_stable = w362;
	assign DRV_LOW_a[10] = w287;
	assign n_DRV_HIGH_a[10] = w34;
	assign w211 = n_INPUT_a[10];
	assign w356 = int_serial;
	assign test_2 = w213;
	assign n_test_reset = w54;
	assign lfo_16384Hz = w53;
	assign sc_write = w315;
	assign w158 = n_INPUT_nrd;
	assign sc_read = w145;
	assign n_DRV_HIGH_nrd = w35;
	assign sb_read = w144;
	assign w74 = clk9;
	assign n_ext_addr_en = w8;
	assign DRV_LOW_nwr = w214;
	assign w215 = n_INPUT_nwr;
	assign DRV_LOW_nrd = w41;
	assign n_DRV_HIGH_nwr = w40;
	assign n_sb_write = w357;
	assign w39 = n_t1_frompad;
	assign w52 = n_t2_frompad;
	assign w63 = n_reset2;
	assign addr_latch = w129;
	assign w85 = int_jp;
	assign w86 = FF60_D1;
	assign test_1 = w36;
	assign dma_addr_ext = w88;
	assign w310 = clk4;
	assign lfo_512Hz = w112;
	assign a[0] = w111;
	assign soc_wr = w109;
	assign a[1] = w107;
	assign a[3] = w247;
	assign a[5] = w106;
	assign a[6] = w248;
	assign a[2] = w304;
	assign a[7] = w249;
	assign a[4] = w102;
	assign d[1] = w68;
	assign d[2] = w71;
	assign d[0] = w31;
	assign d[6] = w117;
	assign d[5] = w19;
	assign d[3] = w23;
	assign d[4] = w94;
	assign d[7] = w153;
	assign soc_rd = w45;
	assign CONST0 = w20;
	assign dma_a[5] = w279;
	assign dma_a[1] = w171;
	assign dma_a[6] = w170;
	assign dma_a[3] = w341;
	assign n_cpu_m1 = w285;
	assign dma_a[2] = w245;
	assign w147 = ffxx;
	assign dma_a[0] = w172;
	assign dma_a[4] = w173;
	assign oam_dma_wr = w342;
	assign dma_a[10] = w280;
	assign dma_a[7] = w177;
	assign w178 = ppu_clk;
	assign w204 = clk6;
	assign dma_a[11] = w205;
	assign w239 = ppu_wr;
	assign w182 = clk6_delay;
	assign dma_a[12] = w156;
	assign dma_run = w183;
	assign w238 = ff46;
	assign dma_a[8] = w237;
	assign n_dma_phi = w321;
	assign w186 = n_ppu_hard_reset;
	assign dma_a[9] = w274;
	assign w284 = cpu_m1;
	assign cpu_vram_oam_rd = w180;
	assign cpu_irq_trig[4] = w130;
	assign w257 = ppu_int_stat;
	assign w131 = cpu_irq_ack[4];
	assign a[10] = w318;
	assign w258 = clk2;
	assign w166 = cpu_irq_ack[3];
	assign vram_to_oam = w167;
	assign w65 = ppu_int_vbl;
	assign w255 = cpu_irq_ack[2];
	assign cpu_irq_trig[1] = w150;
	assign cpu_irq_trig[2] = w151;
	assign cpu_irq_trig[3] = w160;
	assign w161 = cpu_irq_ack[1];
	assign cpu_irq_trig[0] = w162;
	assign w322 = cpu_irq_ack[0];
	assign w261 = non_vram_mreq;
	assign dma_a_15 = w190;
	assign w200 = osc_ena;
	assign a[13] = w4;
	assign w199 = cpu_wr;
	assign n_extdb_to_intdb = w300;
	assign n_dblatch_to_intdb = w260;
	assign w55 = reset;
	assign n_intdb_to_extdb = w259;
	assign w201 = cpu_wr_sync;
	assign a[14] = w28;
	assign n_ena_pu_db = w297;
	assign a[11] = w48;
	assign w47 = cpu_rd;
	assign a[8] = w270;
	assign a[9] = w227;
	assign a[12] = w49;
	assign w293 = n_INPUT_a[12];

	// Instances

	dmg_not g1 (.a(w6), .x(w5) );
	dmg_not g2 (.a(w293), .x(w50) );
	dmg_not g3 (.a(w273), .x(w272) );
	dmg_not g4 (.a(w198), .x(w197) );
	dmg_not g5 (.a(w261), .x(w323) );
	dmg_not g6 (.a(w322), .x(w191) );
	dmg_not g7 (.a(w259), .x(w297) );
	dmg_not g8 (.a(w190), .x(w189) );
	dmg_not g9 (.a(w161), .x(w66) );
	dmg_not g10 (.a(w168), .x(w167) );
	dmg_not g11 (.a(w255), .x(w254) );
	dmg_not g12 (.a(w166), .x(w165) );
	dmg_not g13 (.a(w131), .x(w70) );
	dmg_not g14 (.a(w283), .x(w175) );
	dmg_not g15 (.a(w188), .x(w282) );
	dmg_not g16 (.a(w281), .x(w88) );
	dmg_not g17 (.a(w240), .x(w241) );
	dmg_not g18 (.a(w284), .x(w285) );
	dmg_not g19 (.a(w308), .x(w307) );
	dmg_not g20 (.a(w339), .x(w340) );
	dmg_not g21 (.a(w267), .x(w11) );
	dmg_not g22 (.a(w115), .x(w116) );
	dmg_not g23 (.a(w32), .x(w69) );
	dmg_not g24 (.a(w45), .x(w44) );
	dmg_not g25 (.a(w136), .x(w137) );
	dmg_not g26 (.a(w36), .x(w8) );
	dmg_not g27 (.a(w140), .x(w139) );
	dmg_not g28 (.a(w39), .x(w38) );
	dmg_not g29 (.a(w52), .x(w159) );
	dmg_not g30 (.a(w217), .x(w53) );
	dmg_not g31 (.a(w200), .x(w56) );
	dmg_not g32 (.a(w142), .x(w143) );
	dmg_not g33 (.a(w78), .x(w77) );
	dmg_not g34 (.a(w80), .x(w81) );
	dmg_not g35 (.a(w312), .x(w311) );
	dmg_not g36 (.a(w113), .x(w112) );
	dmg_not g37 (.a(w104), .x(w105) );
	dmg_not g38 (.a(w304), .x(w303) );
	dmg_not g39 (.a(w313), .x(w343) );
	dmg_not g40 (.a(w211), .x(w210) );
	dmg_not g41 (.a(w263), .x(w264) );
	dmg_not g42 (.a(w149), .x(w317) );
	dmg_not g43 (.a(w241), .x(w154) );
	dmg_not g44 (.a(w307), .x(w306) );
	dmg_not g45 (.a(w272), .x(w129) );
	dmg_not g46 (.a(w213), .x(w271) );
	dmg_not g47 (.a(w201), .x(w202) );
	dmg_not g48 (.a(w203), .x(w269) );
	dmg_not g49 (.a(w63), .x(w29) );
	dmg_not g50 (.a(w16), .x(w12) );
	dmg_not g51 (.a(w233), .x(w232) );
	dmg_not g52 (.a(w10), .x(w9) );
	dmg_nor g53 (.a(w36), .b(w2), .x(w1) );
	dmg_nor g54 (.a(w36), .b(w363), .x(w290) );
	dmg_nor g55 (.a(w36), .b(w228), .x(w289) );
	dmg_nor g56 (.a(w258), .b(w36), .x(w344) );
	dmg_nor g57 (.a(w240), .b(w275), .x(w276) );
	dmg_nor g58 (.a(w277), .b(w185), .x(w184) );
	dmg_nor g59 (.a(w29), .b(w354), .x(w15) );
	dmg_nor g60 (.a(w29), .b(w230), .x(w231) );
	dmg_nor g61 (.a(w29), .b(w18), .x(w17) );
	dmg_nor g62 (.a(w29), .b(w90), .x(w91) );
	dmg_nor g63 (.a(w29), .b(w333), .x(w332) );
	dmg_nor g64 (.a(w36), .b(w286), .x(w287) );
	dmg_nor g65 (.a(w88), .b(w43), .x(w42) );
	dmg_nor g66 (.a(w36), .b(w194), .x(w214) );
	dmg_nor g67 (.a(w36), .b(w42), .x(w41) );
	dmg_nor g68 (.a(w132), .b(w126), .x(w125) );
	dmg_nor g69 (.a(w36), .b(w26), .x(w266) );
	dmg_nor g70 (.a(w29), .b(w121), .x(w349) );
	dmg_nor g71 (.a(w29), .b(w120), .x(w348) );
	dmg_nor g72 (.a(w29), .b(w30), .x(w326) );
	dmg_nor g73 (.a(w261), .b(w213), .x(w196) );
	dmg_nor g74 (.a(w14), .b(w13), .x(w355) );
	dmg_nor g75 (.a(w36), .b(w225), .x(w268) );
	dmg_nor g76 (.a(w36), .b(w235), .x(w292) );
	dmg_nand g77 (.a(w2), .b(w8), .x(w7) );
	dmg_nand g78 (.a(w363), .b(w8), .x(w288) );
	dmg_nand g79 (.a(w228), .b(w8), .x(w51) );
	dmg_nand g80 (.a(w36), .b(w259), .x(w300) );
	dmg_nand g81 (.a(w319), .b(w320), .x(w181) );
	dmg_nand g82 (.a(w320), .b(w186), .x(w283) );
	dmg_nand g83 (.a(w194), .b(w8), .x(w40) );
	dmg_nand g84 (.a(w42), .b(w8), .x(w35) );
	dmg_nand g85 (.a(w26), .b(w8), .x(w265) );
	dmg_nand g86 (.a(w309), .b(w182), .x(w179) );
	dmg_nand g87 (.a(w183), .b(w282), .x(w281) );
	dmg_nand g88 (.a(w183), .b(w188), .x(w168) );
	dmg_nand g89 (.a(w225), .b(w8), .x(w234) );
	dmg_nand g90 (.a(w235), .b(w8), .x(w291) );
	dmg_bufif0 g91 (.a0(w50), .n_ena(w8), .a1(w50), .x(w49) );
	dmg_bufif0 g92 (.a0(w5), .n_ena(w8), .a1(w5), .x(w4) );
	dmg_bufif0 g93 (.a0(w232), .n_ena(w8), .a1(w232), .x(w270) );
	dmg_bufif0 g94 (.a0(w9), .n_ena(w8), .a1(w9), .x(w48) );
	dmg_bufif0 g95 (.a0(w11), .n_ena(w8), .a1(w11), .x(w227) );
	dmg_bufif0 g96 (.a0(w264), .n_ena(w8), .a1(w264), .x(w28) );
	dmg_latch g97 (.ena(w129), .d(w49), .q(w207) );
	dmg_latch g98 (.ena(w129), .d(w48), .q(w206) );
	dmg_latch g99 (.ena(w129), .d(w270), .q(w236) );
	dmg_latch g100 (.ena(w129), .d(w4), .q(w3) );
	dmg_latch g101 (.ena(w129), .d(w227), .q(w226) );
	dmg_latch g102 (.ena(w149), .d(w130), .nq(w152) );
	dmg_latch g103 (.ena(w149), .d(w160), .nq(w163) );
	dmg_latch g104 (.ena(w129), .d(w28), .q(w27) );
	dmg_latch g105 (.ena(w149), .d(w150), .nq(w351) );
	dmg_latch g106 (.ena(w149), .d(w162), .nq(w316) );
	dmg_latch g107 (.ena(w129), .d(w318), .q(w337) );
	dmg_latch g108 (.ena(w149), .d(w151), .nq(w324) );
	dmg_bufif0 g109 (.a0(w210), .n_ena(w8), .a1(w210), .x(w318) );
	dmg_dffr g110 (.clk(w74), .nr1(w12), .d(w14), .nr2(w12), .nq(w13) );
	dmg_dffr g111 (.clk(w223), .nr1(w63), .d(w68), .nr2(w63), .nq(w336), .q(w335) );
	dmg_dffr g112 (.clk(w358), .nr1(w175), .d(w169), .nr2(w175), .nq(w169), .q(w170) );
	dmg_dffr g113 (.clk(w365), .nr1(w175), .d(w174), .nr2(w175), .nq(w174), .q(w173) );
	dmg_dffr g114 (.clk(w338), .nr1(w175), .d(w244), .nr2(w175), .nq(w244), .q(w245) );
	dmg_dffr g115 (.clk(w359), .nr1(w175), .d(w278), .nr2(w175), .nq(w278), .q(w172) );
	dmg_dffr g116 (.clk(w277), .nr1(w186), .d(w276), .nr2(w186), .q(w364) );
	dmg_dffr g117 (.clk(w321), .nr1(w186), .d(w364), .nr2(w186), .nq(w320) );
	dmg_dffr g118 (.clk(w79), .nr1(w61), .d(w76), .nr2(w61), .nq(w76), .q(w312) );
	dmg_dffr g119 (.clk(w103), .nr1(w61), .d(w79), .nr2(w61), .nq(w79), .q(w78) );
	dmg_dffr g120 (.clk(w76), .nr1(w61), .d(w314), .nr2(w61), .nq(w314), .q(w313) );
	dmg_dffr g121 (.clk(w314), .nr1(w61), .d(w114), .nr2(w61), .nq(w114), .q(w113) );
	dmg_dffr g122 (.clk(w216), .nr1(w61), .d(w141), .nr2(w61), .nq(w141), .q(w142) );
	dmg_dffr g123 (.clk(w193), .nr1(w61), .d(w75), .nr2(w61), .nq(w75), .q(w217) );
	dmg_dffr g124 (.clk(w223), .nr1(w63), .d(w94), .nr2(w63), .nq(w96), .q(w95) );
	dmg_dffr g125 (.clk(w221), .nr1(w61), .d(w62), .nr2(w61), .nq(w62), .q(w140) );
	dmg_dffr g126 (.clk(w223), .nr1(w63), .d(w23), .nr2(w63), .nq(w329), .q(w222) );
	dmg_dffr g127 (.clk(w328), .nr1(w61), .d(w60), .nr2(w61), .nq(w60), .q(w59) );
	dmg_dffr g128 (.clk(w62), .nr1(w61), .d(w328), .nr2(w61), .nq(w328) );
	dmg_dffr g129 (.clk(w141), .nr1(w61), .d(w193), .nr2(w61), .nq(w193) );
	dmg_dffr g130 (.clk(w37), .nr1(w61), .d(w216), .nr2(w61), .nq(w216) );
	dmg_dffr g131 (.clk(w74), .nr1(w61), .d(w352), .nr2(w61), .nq(w352) );
	dmg_dffr g132 (.clk(w352), .nr1(w61), .d(w37), .nr2(w61), .nq(w37), .q(w80) );
	dmg_dffr g133 (.clk(w87), .nr1(w61), .d(w103), .nr2(w61), .nq(w103), .q(w104) );
	dmg_dffr g134 (.clk(w148), .nr1(w63), .d(w71), .nr2(w63), .nq(w126) );
	dmg_dffr g135 (.clk(w148), .nr1(w63), .d(w31), .nr2(w63), .nq(w345), .q(w82) );
	dmg_dffr g136 (.clk(w148), .nr1(w63), .d(w68), .nr2(w63), .nq(w251), .q(w250) );
	dmg_dffr g137 (.clk(w114), .nr1(w61), .d(w224), .nr2(w61), .nq(w224), .q(w136) );
	dmg_dffr g138 (.clk(w224), .nr1(w61), .d(w221), .nr2(w61), .nq(w221), .q(w115) );
	dmg_dffr g139 (.clk(w223), .nr1(w63), .d(w153), .nr2(w63), .nq(w301), .q(w361) );
	dmg_dffr g140 (.clk(w223), .nr1(w63), .d(w31), .nr2(w63), .nq(w220), .q(w334) );
	dmg_dffr g141 (.clk(w223), .nr1(w63), .d(w19), .nr2(w63), .nq(w97), .q(w98) );
	dmg_dffr g142 (.clk(w223), .nr1(w63), .d(w117), .nr2(w63), .nq(w118), .q(w119) );
	dmg_dffr g143 (.clk(w174), .nr1(w175), .d(w358), .nr2(w175), .nq(w358), .q(w279) );
	dmg_dffr g144 (.clk(w278), .nr1(w175), .d(w338), .nr2(w175), .nq(w338), .q(w171) );
	dmg_dffr g145 (.clk(w178), .nr1(w186), .d(w182), .nr2(w186), .q(w185) );
	dmg_dffr g146 (.clk(w277), .nr1(w186), .d(w181), .nr2(w186), .q(w183) );
	dmg_dffr g147 (.clk(w321), .nr1(w175), .d(w340), .nr2(w175), .nq(w187) );
	dmg_dffr g148 (.clk(w244), .nr1(w175), .d(w365), .nr2(w175), .nq(w365), .q(w341) );
	dmg_dffr g149 (.clk(w169), .nr1(w175), .d(w176), .nr2(w175), .nq(w176), .q(w177) );
	dmg_dffr g150 (.clk(w223), .nr1(w63), .d(w71), .nr2(w63), .nq(w295), .q(w296) );
	dmg_dffr g151 (.clk(w74), .nr1(w63), .d(w355), .nr2(w63), .q(w203) );
	dmg_dffsr g152 (.nset1(w299), .clk(w65), .nres(w64), .q(w162), .nset2(w299), .d(w21) );
	dmg_dffsr g153 (.nset1(w243), .clk(w257), .nres(w256), .q(w150), .nset2(w243), .d(w21) );
	dmg_dffsr g154 (.nset1(w253), .clk(w203), .nres(w350), .q(w151), .nset2(w253), .d(w21) );
	dmg_dffsr g155 (.nset1(w22), .clk(w356), .nres(w192), .q(w160), .nset2(w22), .d(w21) );
	dmg_dffsr g156 (.nset1(w133), .clk(w85), .nres(w134), .q(w130), .nset2(w133), .d(w21) );
	dmg_latchnq_comp g157 (.n_ena(w241), .d(w94), .ena(w154), .q(w156), .nq(w155) );
	dmg_latchnq_comp g158 (.n_ena(w241), .d(w23), .ena(w154), .q(w205), .nq(w353) );
	dmg_latchnq_comp g159 (.n_ena(w241), .d(w31), .ena(w154), .q(w237), .nq(w347) );
	dmg_latchnq_comp g160 (.n_ena(w241), .d(w117), .ena(w154), .q(w325), .nq(w346) );
	dmg_latchnq_comp g161 (.n_ena(w241), .d(w19), .ena(w154), .q(w209), .nq(w252) );
	dmg_latchnq_comp g162 (.n_ena(w241), .d(w68), .ena(w154), .q(w274), .nq(w128) );
	dmg_latchnq_comp g163 (.n_ena(w241), .d(w71), .ena(w154), .q(w280), .nq(w305) );
	dmg_latchnq_comp g164 (.n_ena(w241), .d(w153), .ena(w154), .q(w190), .nq(w242) );
	dmg_aon g165 (.a0(w271), .a1(w261), .b(w213), .x(w273) );
	dmg_aon g166 (.a0(w47), .a1(w323), .b(w199), .x(w198) );
	dmg_cnt g167 (.q(w14), .d(w348), .load(w16), .clk(w123), .nq(w122) );
	dmg_cnt g168 (.q(w124), .d(w326), .load(w16), .clk(w125), .nq(w218) );
	dmg_cnt g169 (.q(w331), .d(w332), .load(w16), .clk(w92), .nq(w93) );
	dmg_cnt g170 (.q(w327), .d(w17), .load(w16), .clk(w331), .nq(w330) );
	dmg_cnt g171 (.q(w92), .d(w91), .load(w16), .clk(w25), .nq(w24) );
	dmg_cnt g172 (.q(w123), .d(w349), .load(w16), .clk(w327), .nq(w229) );
	dmg_cnt g173 (.q(w73), .d(w15), .load(w16), .clk(w124), .nq(w294) );
	dmg_cnt g174 (.q(w25), .d(w231), .load(w16), .clk(w73), .nq(w72) );
	dmg_nor_latch g175 (.s(w240), .r(w283), .nq(w275) );
	dmg_nor_latch g176 (.s(w262), .r(w57), .nq(w58) );
	dmg_muxi g177 (.sel(w99), .d1(w296), .d0(w71), .q(w230) );
	dmg_muxi g178 (.sel(w99), .d1(w361), .d0(w153), .q(w120) );
	dmg_muxi g179 (.sel(w99), .d1(w119), .d0(w117), .q(w121) );
	dmg_muxi g180 (.sel(w99), .d1(w334), .d0(w31), .q(w30) );
	dmg_muxi g181 (.sel(w250), .d1(w83), .d0(w84), .q(w132) );
	dmg_muxi g182 (.sel(w82), .d1(w81), .d0(w77), .q(w84) );
	dmg_muxi g183 (.sel(w82), .d1(w53), .d0(w143), .q(w83) );
	dmg_muxi g184 (.sel(w36), .d1(w158), .d0(w47), .q(w46) );
	dmg_muxi g185 (.sel(w36), .d1(w215), .d0(w201), .q(w157) );
	dmg_muxi g186 (.sel(w99), .d1(w98), .d0(w19), .q(w18) );
	dmg_muxi g187 (.sel(w99), .d1(w222), .d0(w23), .q(w90) );
	dmg_muxi g188 (.sel(w99), .d1(w95), .d0(w94), .q(w333) );
	dmg_muxi g189 (.sel(w99), .d1(w335), .d0(w68), .q(w354) );
	dmg_and g190 (.a(w239), .b(w238), .x(w240) );
	dmg_and g191 (.a(w52), .b(w38), .x(w36) );
	dmg_and g192 (.a(w39), .b(w159), .x(w213) );
	dmg_and g193 (.a(w58), .b(w59), .x(w212) );
	dmg_and g194 (.a(w183), .b(w184), .x(w342) );
	dmg_and g195 (.a(w277), .b(w181), .x(w359) );
	dmg_and g196 (.a(w238), .b(w309), .x(w308) );
	dmg_not2 g197 (.a(w179), .x(w180) );
	dmg_not2 g198 (.a(w277), .x(w321) );
	dmg_not2 g199 (.a(w310), .x(w277) );
	dmg_not g200 (.a(w107), .x(w108) );
	dmg_not g201 (.a(w111), .x(w110) );
	dmg_not3 g202 (.a(w157), .x(w109) );
	dmg_not3 g203 (.a(w46), .x(w45) );
	dmg_and3 g204 (.a(w135), .b(w70), .c(w63), .x(w134) );
	dmg_and4 g205 (.a(w100), .b(w45), .c(w108), .d(w111), .x(w33) );
	dmg_and4 g206 (.a(w100), .b(w45), .c(w107), .d(w110), .x(w89) );
	dmg_and4 g207 (.a(w100), .b(w109), .c(w108), .d(w110), .x(w360) );
	dmg_and4 g208 (.a(w100), .b(w45), .c(w108), .d(w110), .x(w138) );
	dmg_and3 g209 (.a(w164), .b(w165), .c(w63), .x(w192) );
	dmg_and3 g210 (.a(w36), .b(w213), .c(w212), .x(w362) );
	dmg_and4 g211 (.a(w146), .b(w45), .c(w107), .d(w110), .x(w145) );
	dmg_and4 g212 (.a(w146), .b(w45), .c(w108), .d(w111), .x(w144) );
	dmg_notif1 g213 (.ena(w138), .a(w105), .x(w31) );
	dmg_notif1 g214 (.ena(w138), .a(w311), .x(w71) );
	dmg_notif1 g215 (.ena(w138), .a(w343), .x(w23) );
	dmg_notif1 g216 (.ena(w138), .a(w77), .x(w68) );
	dmg_notif1 g217 (.ena(w138), .a(w139), .x(w153) );
	dmg_notif1 g218 (.ena(w33), .a(w72), .x(w71) );
	dmg_notif1 g219 (.ena(w33), .a(w294), .x(w68) );
	dmg_notif1 g220 (.ena(w33), .a(w229), .x(w117) );
	dmg_notif1 g221 (.ena(w89), .a(w118), .x(w117) );
	dmg_notif1 g222 (.ena(w317), .a(w324), .x(w71) );
	dmg_notif1 g223 (.ena(w306), .a(w346), .x(w117) );
	dmg_notif1 g224 (.ena(w306), .a(w252), .x(w19) );
	dmg_notif1 g225 (.ena(w127), .a(w251), .x(w68) );
	dmg_notif1 g226 (.ena(w306), .a(w128), .x(w68) );
	dmg_notif1 g227 (.ena(w127), .a(w345), .x(w31) );
	dmg_notif1 g228 (.ena(w344), .a(w20), .x(w153) );
	dmg_notif1 g229 (.ena(w344), .a(w20), .x(w19) );
	dmg_notif1 g230 (.ena(w344), .a(w20), .x(w117) );
	dmg_notif1 g231 (.ena(w344), .a(w20), .x(w68) );
	dmg_notif1 g232 (.ena(w344), .a(w20), .x(w23) );
	dmg_notif1 g233 (.ena(w344), .a(w20), .x(w71) );
	dmg_notif1 g234 (.ena(w100), .a(w20), .x(w94) );
	dmg_notif1 g235 (.ena(w100), .a(w20), .x(w31) );
	dmg_notif1 g236 (.ena(w306), .a(w305), .x(w71) );
	dmg_notif1 g237 (.ena(w306), .a(w242), .x(w153) );
	dmg_notif1 g238 (.ena(w317), .a(w316), .x(w31) );
	dmg_notif1 g239 (.ena(w317), .a(w351), .x(w68) );
	dmg_notif1 g240 (.ena(w89), .a(w295), .x(w71) );
	dmg_notif1 g241 (.ena(w33), .a(w122), .x(w153) );
	dmg_notif1 g242 (.ena(w89), .a(w336), .x(w68) );
	dmg_notif1 g243 (.ena(w317), .a(w163), .x(w23) );
	dmg_notif1 g244 (.ena(w317), .a(w152), .x(w94) );
	dmg_notif1 g245 (.ena(w306), .a(w347), .x(w31) );
	dmg_notif1 g246 (.ena(w306), .a(w353), .x(w23) );
	dmg_notif1 g247 (.ena(w306), .a(w155), .x(w94) );
	dmg_notif1 g248 (.ena(w127), .a(w126), .x(w71) );
	dmg_notif1 g249 (.ena(w138), .a(w137), .x(w19) );
	dmg_notif1 g250 (.ena(w138), .a(w116), .x(w117) );
	dmg_notif1 g251 (.ena(w89), .a(w301), .x(w153) );
	dmg_notif1 g252 (.ena(w33), .a(w218), .x(w31) );
	dmg_notif1 g253 (.ena(w89), .a(w220), .x(w31) );
	dmg_notif1 g254 (.ena(w33), .a(w93), .x(w94) );
	dmg_notif1 g255 (.ena(w89), .a(w96), .x(w94) );
	dmg_notif1 g256 (.ena(w89), .a(w97), .x(w19) );
	dmg_notif1 g257 (.ena(w33), .a(w330), .x(w19) );
	dmg_notif1 g258 (.ena(w89), .a(w329), .x(w23) );
	dmg_notif1 g259 (.ena(w33), .a(w24), .x(w23) );
	dmg_notif1 g260 (.ena(w138), .a(w112), .x(w94) );
	dmg_nand6 g261 (.a(w172), .b(w171), .c(w245), .d(w341), .e(w173), .f(w177), .x(w339) );
	dmg_nand4 g262 (.a(w101), .b(w246), .c(w147), .d(w45), .x(w149) );
	dmg_nand4 g263 (.a(w101), .b(w246), .c(w147), .d(w109), .x(w32) );
	dmg_mux g264 (.sel(w36), .d1(w44), .d0(w43), .q(w259) );
	dmg_mux g265 (.sel(w86), .d1(w74), .d0(w75), .q(w87) );
	dmg_mux g266 (.sel(w88), .d1(w280), .d0(w337), .q(w286) );
	dmg_mux g267 (.sel(w88), .d1(w325), .d0(w27), .q(w26) );
	dmg_mux g268 (.sel(w88), .d1(w156), .d0(w207), .q(w228) );
	dmg_mux g269 (.sel(w88), .d1(w205), .d0(w206), .q(w363) );
	dmg_mux g270 (.sel(w88), .d1(w237), .d0(w236), .q(w235) );
	dmg_mux g271 (.sel(w88), .d1(w209), .d0(w3), .q(w2) );
	dmg_mux g272 (.sel(w88), .d1(w274), .d0(w226), .q(w225) );
	dmg_nand3 g273 (.a(w181), .b(w187), .c(w186), .x(w319) );
	dmg_nand3 g274 (.a(w47), .b(w261), .c(w204), .x(w260) );
	dmg_and3 g275 (.a(w298), .b(w191), .c(w63), .x(w64) );
	dmg_or g276 (.a(w202), .b(w196), .x(w195) );
	dmg_or g277 (.a(w68), .b(w32), .x(w67) );
	dmg_and3 g278 (.a(w304), .b(w302), .c(w147), .x(w100) );
	dmg_nand g279 (.a(w286), .b(w8), .x(w34) );
	dmg_or g280 (.a(w71), .b(w32), .x(w219) );
	dmg_nand3 g281 (.a(w69), .b(w165), .c(w23), .x(w22) );
	dmg_nand4 g282 (.a(w111), .b(w108), .c(w109), .d(w100), .x(w99) );
	dmg_nand4 g283 (.a(w110), .b(w107), .c(w109), .d(w100), .x(w223) );
	dmg_nand3 g284 (.a(w69), .b(w70), .c(w94), .x(w133) );
	dmg_nand3 g285 (.a(w38), .b(w159), .c(w55), .x(w54) );
	dmg_const g286 (.q0(w20), .q1(w21) );
	dmg_nand3 g287 (.a(w69), .b(w66), .c(w68), .x(w243) );
	dmg_nand3 g288 (.a(w69), .b(w191), .c(w31), .x(w299) );
	dmg_nand3 g289 (.a(w208), .b(w63), .c(w269), .x(w16) );
	dmg_or g290 (.a(w204), .b(w99), .x(w208) );
	dmg_or g291 (.a(w196), .b(w197), .x(w43) );
	dmg_or g292 (.a(w31), .b(w32), .x(w298) );
	dmg_or g293 (.a(w195), .b(w88), .x(w194) );
	dmg_or g294 (.a(w23), .b(w32), .x(w164) );
	dmg_or g295 (.a(w94), .b(w32), .x(w135) );
	dmg_or g296 (.a(w55), .b(w56), .x(w57) );
	dmg_nor5 g297 (.a(w249), .b(w248), .c(w106), .d(w102), .e(w247), .x(w302) );
	dmg_nor4 g298 (.a(w249), .b(w248), .c(w106), .d(w102), .x(w101) );
	dmg_and3 g299 (.a(w303), .b(w302), .c(w147), .x(w146) );
	dmg_and4 g300 (.a(w111), .b(w107), .c(w304), .d(w247), .x(w246) );
	dmg_and4 g301 (.a(w100), .b(w45), .c(w107), .d(w111), .x(w127) );
	dmg_nand4 g302 (.a(w111), .b(w107), .c(w109), .d(w100), .x(w148) );
	dmg_nand3 g303 (.a(w69), .b(w254), .c(w71), .x(w253) );
	dmg_and3 g304 (.a(w219), .b(w254), .c(w63), .x(w350) );
	dmg_nor3 g305 (.a(w209), .b(w325), .c(w189), .x(w188) );
	dmg_and3 g306 (.a(w67), .b(w66), .c(w63), .x(w256) );
	dmg_nand4 g307 (.a(w111), .b(w108), .c(w109), .d(w146), .x(w357) );
	dmg_nand4 g308 (.a(w110), .b(w107), .c(w109), .d(w146), .x(w315) );
	dmg_nor3 g309 (.a(w56), .b(w55), .c(w360), .x(w61) );
endmodule // MMIO