module BootROM (  a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], from_g1_YULA);

	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	input wire a[15];
	input wire from_g1_YULA;

endmodule // BootROM