module MMIO (  reset, clk2, clk4, osc_stable, clk_ena, osc_ena, clk6, clk9, n_reset2, cpu_wr_sync, cpu_m1, n_cpu_m1, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], cpu_irq_trig[4], cpu_irq_ack[4], cpu_irq_trig[3], cpu_irq_ack[3], cpu_irq_trig[2], cpu_irq_ack[2], cpu_irq_trig[1], cpu_irq_ack[1], cpu_irq_trig[0], cpu_irq_ack[0], cpu_rd, cpu_wr, n_DRV_HIGH_a[14], n_INPUT_a[14], DRV_LOW_a[14], n_DRV_HIGH_a[13], n_INPUT_a[13], DRV_LOW_a[13], n_DRV_HIGH_a[12], n_INPUT_a[12], DRV_LOW_a[12], n_DRV_HIGH_a[11], n_INPUT_a[11], DRV_LOW_a[11], n_DRV_HIGH_a[10], n_INPUT_a[10], DRV_LOW_a[10], n_DRV_HIGH_a[9], n_INPUT_a[9], DRV_LOW_a[9], n_DRV_HIGH_a[8], n_INPUT_a[8], DRV_LOW_a[8], n_DRV_HIGH_nrd, n_INPUT_nrd, DRV_LOW_nrd, n_DRV_HIGH_nwr, n_INPUT_nwr, DRV_LOW_nwr, n_t1_frompad, n_t2_frompad, CONST0, n_ena_pu_db, n_dma_phi, dma_a[0], dma_a[4], dma_a[2], dma_a[6], dma_a[10], dma_a[1], dma_a[5], dma_a[11], dma_a[3], dma_a[7], dma_a[8], dma_a[12], dma_a[9], dma_run, soc_wr, soc_rd, lfo_512Hz, ppu_rd, ppu_wr, int_serial, sc_read, sb_read, sc_write, n_sb_write, lfo_16384Hz, ppu_clk, vram_to_oam, dma_a[15], non_vram_mreq, test_1, test_2, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, n_test_reset, n_ext_addr_en, addr_latch, int_jp, FF60_D1, ffxx, n_ppu_hard_reset, ff46, mmio_unk1, cpu_vram_oam_rd, mmio_unk2, ppu_int_stat, ppu_int_vbl, from_ppu2_CATY);

	input wire reset;
	input wire clk2;
	input wire clk4;
	output wire osc_stable;
	input wire clk_ena;
	input wire osc_ena;
	input wire clk6;
	input wire clk9;
	input wire n_reset2;
	input wire cpu_wr_sync;
	input wire cpu_m1;
	output wire n_cpu_m1;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	output wire cpu_irq_trig[4];
	input wire cpu_irq_ack[4];
	output wire cpu_irq_trig[3];
	input wire cpu_irq_ack[3];
	output wire cpu_irq_trig[2];
	input wire cpu_irq_ack[2];
	output wire cpu_irq_trig[1];
	input wire cpu_irq_ack[1];
	output wire cpu_irq_trig[0];
	input wire cpu_irq_ack[0];
	input wire cpu_rd;
	input wire cpu_wr;
	output wire n_DRV_HIGH_a[14];
	input wire n_INPUT_a[14];
	output wire DRV_LOW_a[14];
	output wire n_DRV_HIGH_a[13];
	input wire n_INPUT_a[13];
	output wire DRV_LOW_a[13];
	output wire n_DRV_HIGH_a[12];
	input wire n_INPUT_a[12];
	output wire DRV_LOW_a[12];
	output wire n_DRV_HIGH_a[11];
	input wire n_INPUT_a[11];
	output wire DRV_LOW_a[11];
	output wire n_DRV_HIGH_a[10];
	input wire n_INPUT_a[10];
	output wire DRV_LOW_a[10];
	output wire n_DRV_HIGH_a[9];
	input wire n_INPUT_a[9];
	output wire DRV_LOW_a[9];
	output wire n_DRV_HIGH_a[8];
	input wire n_INPUT_a[8];
	output wire DRV_LOW_a[8];
	output wire n_DRV_HIGH_nrd;
	input wire n_INPUT_nrd;
	output wire DRV_LOW_nrd;
	output wire n_DRV_HIGH_nwr;
	input wire n_INPUT_nwr;
	output wire DRV_LOW_nwr;
	input wire n_t1_frompad;
	input wire n_t2_frompad;
	input wire CONST0;
	output wire n_ena_pu_db;
	output wire n_dma_phi;
	output wire dma_a[0];
	output wire dma_a[4];
	output wire dma_a[2];
	output wire dma_a[6];
	output wire dma_a[10];
	output wire dma_a[1];
	output wire dma_a[5];
	output wire dma_a[11];
	output wire dma_a[3];
	output wire dma_a[7];
	output wire dma_a[8];
	output wire dma_a[12];
	output wire dma_a[9];
	output wire dma_run;
	output wire soc_wr;
	output wire soc_rd;
	output wire lfo_512Hz;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire int_serial;
	output wire sc_read;
	output wire sb_read;
	output wire sc_write;
	output wire n_sb_write;
	output wire lfo_16384Hz;
	input wire ppu_clk;
	output wire vram_to_oam;
	output wire dma_a[15];
	input wire non_vram_mreq;
	output wire test_1;
	output wire test_2;
	output wire n_extdb_to_intdb;
	output wire n_dblatch_to_intdb;
	output wire n_intdb_to_extdb;
	output wire n_test_reset;
	output wire n_ext_addr_en;
	output wire addr_latch;
	input wire int_jp;
	input wire FF60_D1;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ff46;
	output wire mmio_unk1;
	output wire cpu_vram_oam_rd;
	output wire mmio_unk2;
	input wire ppu_int_stat;
	input wire ppu_int_vbl;
	input wire from_ppu2_CATY;

endmodule // MMIO