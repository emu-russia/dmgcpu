module APU (  cclk, clk2, clk4, clk6, clk7, clk9, n_reset2, a, d, cpu_wakeup, n_DRV_HIGH_a, n_INPUT_a, DRV_LOW_a,  
	n_sout_topad, n_DRV_HIGH_sin, n_ENA_PU_sin, DRV_LOW_sin, n_DRV_HIGH_sck, sck_dir, DRV_LOW_sck, n_DRV_HIGH_p10, CONST0, n_p10, DRV_LOW_p10, n_DRV_HIGH_p11, n_p11, DRV_LOW_p11, n_DRV_HIGH_p12, n_p12, DRV_LOW_p12, n_DRV_HIGH_p13, n_p13, DRV_LOW_p13, n_DRV_HIGH_p14, DRV_LOW_p14, n_DRV_HIGH_p15, DRV_LOW_p15, 
	dma_a, soc_wr, soc_rd, lfo_512Hz, ser_out, serial_tick, test_1, test_2, n_ext_addr_en, ch3_active, 
	wave_a, wave_rd, n_wave_wr, wave_bl_pch, n_wave_rd, addr_latch, int_jp, FF60_D1, ffxx, n_ch1_amp_en, n_ch2_amp_en, n_ch3_amp_en, n_ch4_amp_en, 
	ch1_out, ch2_out, ch3_out, ch4_out, r_vin_en, rmixer, l_vin_en, lmixer, n_rvolume, n_lvolume, dma_addr_ext);

	input wire cclk;
	input wire clk2;
	input wire clk4;
	input wire clk6;
	input wire clk7;
	input wire clk9;
	input wire n_reset2;
	inout wire [7:0] a; 			// 7:0 are used only   ⚠️ bidir
	inout wire [7:0] d;
	output wire cpu_wakeup;
	output wire [7:0] n_DRV_HIGH_a;
	input wire [7:0] n_INPUT_a;
	output wire [7:0] DRV_LOW_a;
	output wire n_sout_topad;
	output wire n_DRV_HIGH_sin;
	output wire n_ENA_PU_sin;
	output wire DRV_LOW_sin;
	output wire n_DRV_HIGH_sck;
	input wire sck_dir;
	output wire DRV_LOW_sck;
	output wire n_DRV_HIGH_p10;
	inout wire CONST0;
	input wire n_p10;
	output wire DRV_LOW_p10;
	output wire n_DRV_HIGH_p11;
	input wire n_p11;
	output wire DRV_LOW_p11;
	output wire n_DRV_HIGH_p12;
	input wire n_p12;
	output wire DRV_LOW_p12;
	output wire n_DRV_HIGH_p13;
	input wire n_p13;
	output wire DRV_LOW_p13;
	output wire n_DRV_HIGH_p14;
	output wire DRV_LOW_p14;
	output wire n_DRV_HIGH_p15;
	output wire DRV_LOW_p15;
	input wire [7:0] dma_a; 		// 7:0 are used only
	input wire soc_wr;
	input wire soc_rd;
	input wire lfo_512Hz;
	input wire ser_out;
	input wire serial_tick;
	input wire test_1;
	input wire test_2;
	input wire n_ext_addr_en;
	output wire ch3_active;
	output wire [3:0] wave_a;
	input wire [7:0] wave_rd;
	output wire n_wave_wr;
	output wire wave_bl_pch;
	output wire n_wave_rd;
	input wire addr_latch;
	output wire int_jp;
	output wire FF60_D1;
	input wire ffxx;
	output wire n_ch1_amp_en;
	output wire n_ch2_amp_en;
	output wire n_ch3_amp_en;
	output wire n_ch4_amp_en;
	output wire [3:0] ch1_out;
	output wire [3:0] ch2_out;
	output wire [3:0] ch3_out;
	output wire [3:0] ch4_out;
	output wire r_vin_en;
	output wire [3:0] rmixer;
	output wire l_vin_en;
	output wire [3:0] lmixer;
	output wire [2:0] n_rvolume;
	output wire [2:0] n_lvolume;
	input wire dma_addr_ext;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire w1083;
	wire w1084;
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;

	assign w1144 = n_INPUT_a[5];
	assign n_DRV_HIGH_a[5] = w1145;
	assign DRV_LOW_a[6] = w1244;
	assign DRV_LOW_a[5] = w2;
	assign w1 = n_INPUT_a[4];
	assign w88 = n_INPUT_a[6];
	assign n_DRV_HIGH_a[6] = w1243;
	assign DRV_LOW_a[7] = w89;
	assign w702 = n_INPUT_a[7];
	assign n_DRV_HIGH_a[4] = w703;
	assign DRV_LOW_a[1] = w621;
	assign DRV_LOW_a[4] = w622;
	assign n_DRV_HIGH_a[3] = w1249;
	assign n_DRV_HIGH_a[7] = w1148;
	assign w1147 = n_INPUT_a[3];
	assign DRV_LOW_a[3] = w661;
	assign n_DRV_HIGH_a[2] = w1039;
	assign w660 = n_INPUT_a[2];
	assign DRV_LOW_a[2] = w1040;
	assign n_DRV_HIGH_a[1] = w701;
	assign w700 = n_INPUT_a[1];
	assign w444 = n_INPUT_a[0];
	assign n_DRV_HIGH_a[0] = w126;
	assign DRV_LOW_a[0] = w127;
	assign n_sout_topad = w1233;
	assign n_DRV_HIGH_sin = w804;
	assign DRV_LOW_sin = w802;
	assign n_DRV_HIGH_sck = w882;
	assign DRV_LOW_sck = w1273;
	assign n_ENA_PU_sin = w618;
	assign n_DRV_HIGH_p10 = w937;
	assign DRV_LOW_p10 = w564;
	assign n_DRV_HIGH_p13 = w939;
	assign n_DRV_HIGH_p11 = w877;
	assign DRV_LOW_p13 = w938;
	assign DRV_LOW_p11 = w561;
	assign n_DRV_HIGH_p14 = w562;
	assign DRV_LOW_p14 = w620;
	assign w777 = n_p10;
	assign n_DRV_HIGH_p12 = w435;
	assign w778 = n_p11;
	assign w780 = n_p13;
	assign DRV_LOW_p12 = w876;
	assign w781 = n_p12;
	assign DRV_LOW_p15 = w797;
	assign n_DRV_HIGH_p15 = w832;
	assign n_lvolume[2] = w224;
	assign n_rvolume[2] = w1153;
	assign n_rvolume[1] = w376;
	assign n_lvolume[1] = w1151;
	assign n_rvolume[0] = w227;
	assign n_lvolume[0] = w226;
	assign l_vin_en = w1109;
	assign ch4_out[3] = w1152;
	assign ch4_out[2] = w131;
	assign ch4_out[1] = w130;
	assign lmixer[1] = w1072;
	assign ch4_out[0] = w1071;
	assign lmixer[0] = w1094;
	assign rmixer[1] = w1108;
	assign r_vin_en = w815;
	assign lmixer[2] = w1047;
	assign rmixer[2] = w816;
	assign lmixer[3] = w1048;
	assign rmixer[3] = w17;
	assign rmixer[0] = w18;
	assign n_ch4_amp_en = w836;
	assign CONST0 = w20;
	assign ch2_out[3] = w1344;
	assign ch2_out[2] = w1345;
	assign ch2_out[1] = w1328;
	assign n_ch1_amp_en = w529;
	assign ch2_out[0] = w1343;
	assign ch1_out[1] = w545;
	assign w1317 = lfo_512Hz;
	assign ch1_out[0] = w544;
	assign ch1_out[2] = w543;
	assign ch1_out[3] = w542;
	assign w114 = soc_rd;
	assign d[3] = w229;
	assign d[6] = w55;
	assign d[5] = w16;
	assign d[2] = w180;
	assign d[7] = w187;
	assign d[0] = w183;
	assign w800 = soc_wr;
	assign w7 = dma_a[0];
	assign w880 = ffxx;
	assign w881 = sck_dir;
	assign w1202 = clk6;
	assign d[4] = w29;
	assign d[1] = w331;
	assign w8 = clk7;
	assign ch3_out[3] = w714;
	assign ch3_out[2] = w1037;
	assign ch3_out[1] = w1334;
	assign cpu_wakeup = w1203;
	assign a[7] = w666;
	assign w559 = n_reset2;
	assign n_ch2_amp_en = w755;
	assign ch3_out[0] = w754;
	assign w57 = ser_out;
	assign a[6] = w112;
	assign a[4] = w111;
	assign n_ch3_amp_en = w408;
	assign a[2] = w104;
	assign a[5] = w578;
	assign w579 = dma_a[4];
	assign w691 = dma_a[2];
	assign a[3] = w110;
	assign w1330 = test_2;
	assign w11 = clk2;
	assign w10 = clk9;
	assign a[1] = w103;
	assign int_jp = w1038;
	assign w383 = dma_addr_ext;
	assign FF60_D1 = w712;
	assign w385 = dma_a[7];
	assign w386 = cclk;
	assign a[0] = w667;
	assign w1126 = serial_tick;
	assign w1125 = dma_a[3];
	assign w1341 = dma_a[5];
	assign w576 = dma_a[6];
	assign w381 = dma_a[1];
	assign w380 = wave_rd[4];
	assign n_wave_wr = w575;
	assign w1157 = wave_rd[5];
	assign w5 = addr_latch;
	assign n_wave_rd = w705;
	assign w583 = wave_rd[7];
	assign w584 = wave_rd[3];
	assign w403 = wave_rd[1];
	assign wave_bl_pch = w1163;
	assign w1162 = wave_rd[6];
	assign w573 = wave_rd[2];
	assign w90 = test_1;
	assign w514 = wave_rd[0];
	assign ch3_active = w397;
	assign w125 = n_ext_addr_en;
	assign wave_a[3] = w1143;
	assign wave_a[2] = w1142;
	assign wave_a[1] = w1340;
	assign wave_a[0] = w1141;
	assign w123 = clk4;

	// Instances

	dmg_not g1 (.a(w1), .x(w124) );
	dmg_not g2 (.a(w388), .x(w960) );
	dmg_not g3 (.a(w388), .x(w961) );
	dmg_not g4 (.a(w1144), .x(w1161) );
	dmg_not g5 (.a(w573), .x(w572) );
	dmg_not g6 (.a(w1158), .x(w708) );
	dmg_not g7 (.a(w70), .x(w519) );
	dmg_not g8 (.a(w388), .x(w1165) );
	dmg_not g9 (.a(w70), .x(w696) );
	dmg_not g10 (.a(w583), .x(w756) );
	dmg_not g11 (.a(w584), .x(w757) );
	dmg_not g12 (.a(w1158), .x(w1159) );
	dmg_not g13 (.a(w704), .x(w706) );
	dmg_not g14 (.a(w386), .x(w387) );
	dmg_not g15 (.a(w70), .x(w40) );
	dmg_not g16 (.a(w957), .x(w1196) );
	dmg_not g17 (.a(w111), .x(w710) );
	dmg_not g18 (.a(w666), .x(w1204) );
	dmg_not g19 (.a(w112), .x(w1200) );
	dmg_not g20 (.a(w11), .x(w12) );
	dmg_not g21 (.a(w8), .x(w580) );
	dmg_not g22 (.a(w112), .x(w113) );
	dmg_not g23 (.a(w931), .x(w932) );
	dmg_not g24 (.a(w70), .x(w942) );
	dmg_not g25 (.a(w70), .x(w1025) );
	dmg_not g26 (.a(w388), .x(w1051) );
	dmg_not g27 (.a(w76), .x(w223) );
	dmg_not g28 (.a(w70), .x(w1106) );
	dmg_not g29 (.a(w69), .x(w1107) );
	dmg_not g30 (.a(w44), .x(w830) );
	dmg_not g31 (.a(w44), .x(w829) );
	dmg_not g32 (.a(w826), .x(w827) );
	dmg_not g33 (.a(w78), .x(w79) );
	dmg_not g34 (.a(w1027), .x(w1028) );
	dmg_not g35 (.a(w1089), .x(w1026) );
	dmg_not g36 (.a(w282), .x(w283) );
	dmg_not g37 (.a(w166), .x(w167) );
	dmg_not g38 (.a(w291), .x(w1316) );
	dmg_not g39 (.a(w144), .x(w299) );
	dmg_not g40 (.a(w144), .x(w930) );
	dmg_not g41 (.a(w44), .x(w1131) );
	dmg_not g42 (.a(w217), .x(w1307) );
	dmg_not g43 (.a(w83), .x(w287) );
	dmg_not g44 (.a(w997), .x(w998) );
	dmg_not g45 (.a(w1305), .x(w1304) );
	dmg_not g46 (.a(w1190), .x(w1189) );
	dmg_not g47 (.a(w167), .x(w168) );
	dmg_not g48 (.a(w943), .x(w992) );
	dmg_not g49 (.a(w70), .x(w946) );
	dmg_not g50 (.a(w1293), .x(w1294) );
	dmg_not g51 (.a(w1006), .x(w1007) );
	dmg_not g52 (.a(w44), .x(w1176) );
	dmg_not g53 (.a(w65), .x(w66) );
	dmg_not g54 (.a(w70), .x(w626) );
	dmg_not g55 (.a(w963), .x(w1302) );
	dmg_not g56 (.a(w493), .x(w1299) );
	dmg_not g57 (.a(w84), .x(w83) );
	dmg_not g58 (.a(w887), .x(w317) );
	dmg_not g59 (.a(w1207), .x(w38) );
	dmg_not g60 (.a(w88), .x(w989) );
	dmg_not g61 (.a(w702), .x(w87) );
	dmg_not g62 (.a(w403), .x(w377) );
	dmg_not g63 (.a(w379), .x(w378) );
	dmg_not g64 (.a(w514), .x(w513) );
	dmg_not g65 (.a(w551), .x(w646) );
	dmg_not g66 (.a(w1162), .x(w645) );
	dmg_not g67 (.a(w70), .x(w1246) );
	dmg_not g68 (.a(w700), .x(w699) );
	dmg_not g69 (.a(w388), .x(w390) );
	dmg_not g70 (.a(w70), .x(w1320) );
	dmg_not g71 (.a(w70), .x(w1319) );
	dmg_not g72 (.a(w388), .x(w389) );
	dmg_not g73 (.a(w744), .x(w745) );
	dmg_not g74 (.a(w1212), .x(w1213) );
	dmg_not g75 (.a(w1241), .x(w1290) );
	dmg_not g76 (.a(w551), .x(w550) );
	dmg_not g77 (.a(w406), .x(w405) );
	dmg_not g78 (.a(w397), .x(w398) );
	dmg_not g79 (.a(w915), .x(w170) );
	dmg_not g80 (.a(w70), .x(w152) );
	dmg_not g81 (.a(w229), .x(w1184) );
	dmg_not g82 (.a(w144), .x(w765) );
	dmg_not g83 (.a(w320), .x(w319) );
	dmg_not g84 (.a(w838), .x(w1367) );
	dmg_not g85 (.a(w42), .x(w43) );
	dmg_not g86 (.a(w821), .x(w1358) );
	dmg_not g87 (.a(w476), .x(w119) );
	dmg_not g88 (.a(w119), .x(w118) );
	dmg_not g89 (.a(w809), .x(w808) );
	dmg_not g90 (.a(w858), .x(w857) );
	dmg_not g91 (.a(w324), .x(w325) );
	dmg_not g92 (.a(w823), .x(w473) );
	dmg_not g93 (.a(w886), .x(w822) );
	dmg_not g94 (.a(w151), .x(w885) );
	dmg_not g95 (.a(w331), .x(w327) );
	dmg_not g96 (.a(w70), .x(w121) );
	dmg_not g97 (.a(w1194), .x(w1193) );
	dmg_not g98 (.a(w70), .x(w1192) );
	dmg_not g99 (.a(w918), .x(w917) );
	dmg_not g100 (.a(w1281), .x(w1280) );
	dmg_not g101 (.a(w915), .x(w916) );
	dmg_not g102 (.a(w537), .x(w538) );
	dmg_not g103 (.a(w915), .x(w1219) );
	dmg_not g104 (.a(w44), .x(w1221) );
	dmg_not g105 (.a(w210), .x(w1220) );
	dmg_not g106 (.a(w44), .x(w500) );
	dmg_not g107 (.a(w1130), .x(w1276) );
	dmg_not g108 (.a(w902), .x(w1253) );
	dmg_not g109 (.a(w44), .x(w400) );
	dmg_not g110 (.a(w504), .x(w721) );
	dmg_not g111 (.a(w501), .x(w1339) );
	dmg_not g112 (.a(w70), .x(w1354) );
	dmg_not g113 (.a(w1355), .x(w1356) );
	dmg_not g114 (.a(w551), .x(w456) );
	dmg_not g115 (.a(w525), .x(w552) );
	dmg_not g116 (.a(w1382), .x(w1383) );
	dmg_not g117 (.a(w556), .x(w555) );
	dmg_not g118 (.a(w679), .x(w680) );
	dmg_not g119 (.a(w598), .x(w738) );
	dmg_not g120 (.a(w70), .x(w594) );
	dmg_not g121 (.a(w70), .x(w600) );
	dmg_not g122 (.a(w1260), .x(w659) );
	dmg_not g123 (.a(w345), .x(w735) );
	dmg_not g124 (.a(w603), .x(w604) );
	dmg_not g125 (.a(w366), .x(w365) );
	dmg_not g126 (.a(w674), .x(w675) );
	dmg_not g127 (.a(w44), .x(w730) );
	dmg_not g128 (.a(w44), .x(w723) );
	dmg_not g129 (.a(w70), .x(w363) );
	dmg_not g130 (.a(w957), .x(w1275) );
	dmg_not g131 (.a(w1223), .x(w1222) );
	dmg_not g132 (.a(w16), .x(w1232) );
	dmg_not g133 (.a(w618), .x(w1231) );
	dmg_not g134 (.a(w881), .x(w1230) );
	dmg_not g135 (.a(w860), .x(w270) );
	dmg_not g136 (.a(w233), .x(w236) );
	dmg_not g137 (.a(w476), .x(w1390) );
	dmg_not g138 (.a(w1011), .x(w1012) );
	dmg_not g139 (.a(w48), .x(w1013) );
	dmg_not g140 (.a(w1013), .x(w1014) );
	dmg_not g141 (.a(w44), .x(w1392) );
	dmg_not g142 (.a(w42), .x(w45) );
	dmg_not g143 (.a(w44), .x(w336) );
	dmg_not g144 (.a(w334), .x(w335) );
	dmg_not g145 (.a(w70), .x(w139) );
	dmg_not g146 (.a(w50), .x(w49) );
	dmg_not g147 (.a(w118), .x(w50) );
	dmg_not g148 (.a(w774), .x(w775) );
	dmg_not g149 (.a(w254), .x(w865) );
	dmg_not g150 (.a(w233), .x(w234) );
	dmg_not g151 (.a(w233), .x(w933) );
	dmg_not g152 (.a(w144), .x(w468) );
	dmg_not g153 (.a(w370), .x(w371) );
	dmg_not g154 (.a(w256), .x(w255) );
	dmg_not g155 (.a(w618), .x(w563) );
	dmg_not g156 (.a(w44), .x(w1335) );
	dmg_not g157 (.a(w1224), .x(w1223) );
	dmg_not g158 (.a(w724), .x(w1227) );
	dmg_not g159 (.a(w70), .x(w1226) );
	dmg_not g160 (.a(w29), .x(w466) );
	dmg_not g161 (.a(w444), .x(w443) );
	dmg_not g162 (.a(w70), .x(w725) );
	dmg_not g163 (.a(w465), .x(w726) );
	dmg_not g164 (.a(w203), .x(w202) );
	dmg_not g165 (.a(w726), .x(w727) );
	dmg_not g166 (.a(w70), .x(w194) );
	dmg_not g167 (.a(w70), .x(w458) );
	dmg_not g168 (.a(w451), .x(w450) );
	dmg_not g169 (.a(w462), .x(w461) );
	dmg_not g170 (.a(w70), .x(w197) );
	dmg_not g171 (.a(w345), .x(w196) );
	dmg_not g172 (.a(w345), .x(w198) );
	dmg_not g173 (.a(w186), .x(w185) );
	dmg_not g174 (.a(w1259), .x(w1260) );
	dmg_not g175 (.a(w602), .x(w601) );
	dmg_not g176 (.a(w181), .x(w182) );
	dmg_not g177 (.a(w70), .x(w749) );
	dmg_not g178 (.a(w452), .x(w906) );
	dmg_not g179 (.a(w70), .x(w430) );
	dmg_not g180 (.a(w957), .x(w958) );
	dmg_not g181 (.a(w70), .x(w1217) );
	dmg_not g182 (.a(w210), .x(w211) );
	dmg_not g183 (.a(w144), .x(w768) );
	dmg_not g184 (.a(w470), .x(w469) );
	dmg_not g185 (.a(w853), .x(w854) );
	dmg_not g186 (.a(w567), .x(w792) );
	dmg_not g187 (.a(w789), .x(w790) );
	dmg_not g188 (.a(w1359), .x(w1360) );
	dmg_not g189 (.a(w70), .x(w52) );
	dmg_not g190 (.a(w136), .x(w137) );
	dmg_not g191 (.a(w70), .x(w338) );
	dmg_not g192 (.a(w320), .x(w72) );
	dmg_not g193 (.a(w44), .x(w820) );
	dmg_not g194 (.a(w70), .x(w262) );
	dmg_not g195 (.a(w219), .x(w218) );
	dmg_not g196 (.a(w874), .x(w873) );
	dmg_not g197 (.a(w161), .x(w845) );
	dmg_not g198 (.a(w409), .x(w410) );
	dmg_not g199 (.a(w1278), .x(w1277) );
	dmg_not g200 (.a(w70), .x(w509) );
	dmg_not g201 (.a(w902), .x(w901) );
	dmg_not g202 (.a(w92), .x(w93) );
	dmg_not g203 (.a(w904), .x(w905) );
	dmg_not g204 (.a(w1251), .x(w548) );
	dmg_not g205 (.a(w180), .x(w527) );
	dmg_not g206 (.a(w638), .x(w1250) );
	dmg_not g207 (.a(w686), .x(w1288) );
	dmg_not g208 (.a(w1261), .x(w684) );
	dmg_not g209 (.a(w659), .x(w746) );
	dmg_not g210 (.a(w100), .x(w101) );
	dmg_not g211 (.a(w405), .x(w404) );
	dmg_not g212 (.a(w1172), .x(w1150) );
	dmg_not g213 (.a(w1290), .x(w1207) );
	dmg_not g214 (.a(w44), .x(w1120) );
	dmg_not g215 (.a(w644), .x(w895) );
	dmg_not g216 (.a(w32), .x(w893) );
	dmg_not g217 (.a(w55), .x(w31) );
	dmg_not g218 (.a(w624), .x(w625) );
	dmg_not g219 (.a(w183), .x(w512) );
	dmg_not g220 (.a(w1175), .x(w1174) );
	dmg_not g221 (.a(w168), .x(w169) );
	dmg_not g222 (.a(w510), .x(w511) );
	dmg_not g223 (.a(w70), .x(w964) );
	dmg_not g224 (.a(w924), .x(w965) );
	dmg_not g225 (.a(w187), .x(w763) );
	dmg_not g226 (.a(w764), .x(w966) );
	dmg_not g227 (.a(w1179), .x(w1180) );
	dmg_not g228 (.a(w161), .x(w160) );
	dmg_not g229 (.a(w912), .x(w910) );
	dmg_not g230 (.a(w161), .x(w913) );
	dmg_not g231 (.a(w320), .x(w321) );
	dmg_not g232 (.a(w969), .x(w968) );
	dmg_not g233 (.a(w286), .x(w285) );
	dmg_not g234 (.a(w219), .x(w280) );
	dmg_not g235 (.a(w833), .x(w615) );
	dmg_not g236 (.a(w839), .x(w838) );
	dmg_not g237 (.a(w986), .x(w987) );
	dmg_not g238 (.a(w70), .x(w1046) );
	dmg_not g239 (.a(w44), .x(w1091) );
	dmg_not g240 (.a(w297), .x(w1044) );
	dmg_not g241 (.a(w313), .x(w312) );
	dmg_not g242 (.a(w1310), .x(w21) );
	dmg_not g243 (.a(w331), .x(w1347) );
	dmg_not g244 (.a(w183), .x(w1348) );
	dmg_not g245 (.a(w282), .x(w281) );
	dmg_not g246 (.a(w115), .x(w116) );
	dmg_not g247 (.a(w44), .x(w1098) );
	dmg_not g248 (.a(w1035), .x(w1097) );
	dmg_not g249 (.a(w886), .x(w1099) );
	dmg_not g250 (.a(w944), .x(w945) );
	dmg_not g251 (.a(w578), .x(w951) );
	dmg_not g252 (.a(w800), .x(w799) );
	dmg_not g253 (.a(w880), .x(w1198) );
	dmg_not g254 (.a(w948), .x(w947) );
	dmg_not g255 (.a(w948), .x(w952) );
	dmg_not g256 (.a(w949), .x(w950) );
	dmg_not g257 (.a(w948), .x(w1264) );
	dmg_not g258 (.a(w1205), .x(w949) );
	dmg_not g259 (.a(w70), .x(w59) );
	dmg_not g260 (.a(w44), .x(w412) );
	dmg_not g261 (.a(w578), .x(w711) );
	dmg_not g262 (.a(w1122), .x(w663) );
	dmg_not g263 (.a(w44), .x(w1121) );
	dmg_not g264 (.a(w1157), .x(w1156) );
	dmg_not g265 (.a(w380), .x(w1155) );
	dmg_not g266 (.a(w1158), .x(w571) );
	dmg_not g267 (.a(w758), .x(w1333) );
	dmg_not g268 (.a(w379), .x(w753) );
	dmg_not g269 (.a(w379), .x(w516) );
	dmg_not g270 (.a(w379), .x(w515) );
	dmg_not g271 (.a(w97), .x(w98) );
	dmg_not g272 (.a(w70), .x(w697) );
	dmg_not g273 (.a(w1147), .x(w689) );
	dmg_not g274 (.a(w660), .x(w1146) );
	dmg_not g275 (.a(w70), .x(w688) );
	dmg_not g276 (.a(w70), .x(w1135) );
	dmg_not g277 (.a(w1137), .x(w1138) );
	dmg_not g278 (.a(w70), .x(w1140) );
	dmg_dffr g279 (.clk(w960), .nr1(w1135), .nr2(w1135), .d(w1136), .q(w1137), .nq(w1136) );
	dmg_dffr g280 (.clk(w961), .nr1(w697), .nr2(w697), .d(w393), .q(w394) );
	dmg_dffr g281 (.clk(w388), .nr2(w697), .d(w392), .q(w393), .nq(w698), .nr1(w697) );
	dmg_dffr g282 (.clk(w1165), .nr1(w696), .nr2(w696), .d(w1166), .q(w282), .nq(w1166) );
	dmg_dffr g283 (.clk(w1196), .nr1(w59), .nr2(w59), .d(w58), .q(w1205), .nq(w58) );
	dmg_dffr g284 (.clk(w1199), .nr1(w559), .nr2(w559), .d(w331), .q(w712) );
	dmg_dffr g285 (.clk(w10), .nr1(w559), .nr2(w559), .d(w9), .q(w713) );
	dmg_dffr g286 (.clk(w10), .nr1(w559), .nr2(w559), .d(w955), .q(w9) );
	dmg_dffr g287 (.clk(w10), .nr1(w559), .nr2(w559), .d(w798), .q(w955) );
	dmg_dffr g288 (.clk(w1051), .nr1(w1046), .nr2(w1046), .d(w1050), .nq(w1050) );
	dmg_dffr g289 (.clk(w1050), .nr1(w1046), .nr2(w1046), .d(w1095), .q(w839), .nq(w1095) );
	dmg_dffr g290 (.clk(w986), .nr1(w818), .nr2(w818), .d(w1112), .q(w1018), .nq(w1112) );
	dmg_dffr g291 (.clk(w284), .nr1(w1025), .nr2(w1025), .d(w1024), .nq(w1024) );
	dmg_dffr g292 (.clk(w1189), .nr1(w164), .nr2(w164), .d(w165), .q(w166), .nq(w165) );
	dmg_dffr g293 (.clk(w570), .nr1(w559), .nr2(w559), .d(w16), .nq(w797) );
	dmg_dffr g294 (.clk(w281), .nr1(w942), .nr2(w942), .d(w295), .nq(w295) );
	dmg_dffr g295 (.clk(w1265), .nr1(w26), .nr2(w26), .d(w25), .q(w24), .nq(w25) );
	dmg_dffr g296 (.clk(w38), .nr1(w40), .nr2(w40), .d(w39), .q(w644), .nq(w39) );
	dmg_dffr g297 (.clk(w1167), .nr1(w1169), .nr2(w1169), .d(w1168), .q(w760), .nq(w1168) );
	dmg_dffr g298 (.clk(w1242), .nr1(w1320), .nr2(w1320), .d(w96), .q(w97) );
	dmg_dffr g299 (.clk(w389), .nr1(w688), .nr2(w688), .d(w687), .q(w686), .nq(w687) );
	dmg_dffr g300 (.clk(w1138), .nr1(w1140), .nr2(w1140), .d(w1139), .q(w1242), .nq(w1139) );
	dmg_dffr g301 (.clk(w1242), .nr1(w744), .nr2(w744), .d(w743), .q(w347) );
	dmg_dffr g302 (.clk(w746), .nr1(w108), .nr2(w108), .d(w1262), .q(w521), .nq(w1262) );
	dmg_dffr g303 (.clk(w1262), .nr1(w108), .nr2(w108), .d(w669), .q(w668), .nq(w669) );
	dmg_dffr g304 (.clk(w669), .nr1(w108), .nr2(w108), .d(w107), .q(w102), .nq(w107) );
	dmg_dffr g305 (.clk(w107), .nr1(w108), .nr2(w108), .d(w106), .q(w105), .nq(w106) );
	dmg_dffr g306 (.clk(w106), .nr1(w108), .nr2(w108), .d(w654), .q(w109), .nq(w654) );
	dmg_dffr g307 (.clk(w169), .nr1(w626), .nr2(w626), .d(w490), .q(w491), .nq(w490) );
	dmg_dffr g308 (.clk(w122), .nr1(w964), .nr2(w964), .d(w922), .q(w920) );
	dmg_dffr g309 (.clk(w149), .nr1(w818), .nr2(w818), .d(w844), .q(w843), .nq(w844) );
	dmg_dffr g310 (.clk(w278), .nr1(w818), .nr2(w818), .d(w279), .q(w1009), .nq(w279) );
	dmg_dffr g311 (.clk(w1058), .nr1(w818), .nr2(w818), .d(w1059), .q(w985), .nq(w1059) );
	dmg_dffr g312 (.clk(w1059), .nr1(w818), .nr2(w818), .d(w1055), .q(w1054), .nq(w1055) );
	dmg_dffr g313 (.clk(w1367), .nr1(w479), .nr2(w479), .d(w1375), .q(w271) );
	dmg_dffr g314 (.clk(w141), .nr1(w262), .nr2(w262), .d(w71), .q(w1359) );
	dmg_dffr g315 (.clk(w141), .nr1(w262), .nr2(w262), .d(w340), .q(w71) );
	dmg_dffr g316 (.clk(w141), .nr1(w853), .nr2(w853), .d(w855), .q(w340) );
	dmg_dffr g317 (.clk(w122), .nr1(w121), .nr2(w121), .d(w260), .q(w120) );
	dmg_dffr g318 (.clk(w1383), .nr1(w671), .nr2(w671), .d(w1353), .q(w1241), .nq(w1353) );
	dmg_dffr g319 (.clk(w1288), .nr1(w598), .nr2(w598), .d(w737), .q(w346) );
	dmg_dffr g320 (.clk(w1288), .nr1(w600), .nr2(w600), .d(w346), .q(w599) );
	dmg_dffr g321 (.clk(w686), .nr1(w600), .nr2(w600), .d(w599), .q(w1261) );
	dmg_dffr g322 (.clk(w367), .nr1(w678), .nr2(w678), .d(w677), .q(w679) );
	dmg_dffr g323 (.clk(w958), .nr1(w725), .nr2(w725), .d(w1236), .q(w465), .nq(w1236) );
	dmg_dffr g324 (.clk(w570), .nr1(w559), .nr2(w559), .d(w183), .q(w846) );
	dmg_dffr g325 (.clk(w570), .nr1(w559), .nr2(w559), .d(w180), .q(w619) );
	dmg_dffr g326 (.clk(w118), .nr1(w242), .nr2(w242), .d(w249), .q(w247) );
	dmg_dffr g327 (.clk(w118), .nr1(w242), .nr2(w242), .d(w246), .q(w249) );
	dmg_dffr g328 (.clk(w118), .nr1(w242), .nr2(w242), .d(w1366), .q(w784) );
	dmg_dffr g329 (.clk(w118), .nr1(w242), .nr2(w242), .d(w1364), .q(w1365) );
	dmg_dffr g330 (.clk(w838), .nr1(w139), .nr2(w139), .d(w140), .q(w1363), .nq(w140) );
	dmg_dffr g331 (.clk(w1390), .nr1(w242), .nr2(w242), .d(w1376), .q(w51) );
	dmg_dffr g332 (.clk(w49), .nr1(w242), .nr2(w242), .d(w51), .q(w243) );
	dmg_dffr g333 (.clk(w49), .nr1(w242), .nr2(w242), .d(w243), .q(w245) );
	dmg_dffr g334 (.clk(w49), .nr1(w242), .nr2(w242), .d(w245), .q(w244) );
	dmg_dffr g335 (.clk(w49), .nr1(w242), .nr2(w242), .d(w244), .q(w241) );
	dmg_dffr g336 (.clk(w49), .nr1(w242), .nr2(w242), .d(w241), .q(w1364) );
	dmg_dffr g337 (.clk(w369), .nr1(w425), .nr2(w425), .d(w424), .q(w565) );
	dmg_dffr g338 (.clk(w367), .nr1(w878), .nr2(w878), .d(w1229), .q(w369) );
	dmg_dffr g339 (.clk(w570), .nr1(w559), .nr2(w559), .d(w331), .q(w560) );
	dmg_dffr g340 (.clk(w570), .nr1(w559), .nr2(w559), .d(w29), .nq(w620) );
	dmg_dffr g341 (.clk(w570), .nr1(w559), .nr2(w559), .d(w187), .q(w803) );
	dmg_dffr g342 (.clk(w570), .nr1(w559), .nr2(w559), .d(w229), .q(w1381) );
	dmg_dffr g343 (.clk(w570), .nr1(w559), .nr2(w559), .d(w55), .q(w56) );
	dmg_dffr g344 (.clk(w1275), .nr1(w1226), .nr2(w1226), .d(w1225), .q(w1224), .nq(w1225) );
	dmg_dffr g345 (.clk(w601), .nr1(w596), .nr2(w596), .d(w1372), .q(w1259), .nq(w1372) );
	dmg_dffr g346 (.clk(w679), .nr1(w95), .nr2(w95), .d(w94), .q(w733) );
	dmg_dffr g347 (.clk(w1255), .nr1(w1276), .nr2(w1276), .d(w187), .nq(w1235) );
	dmg_dffr g348 (.clk(w118), .nr1(w242), .nr2(w242), .d(w1365), .q(w1366) );
	dmg_dffr g349 (.clk(w476), .nr1(w242), .nr2(w242), .d(w247), .q(w248) );
	dmg_dffr g350 (.clk(w476), .nr1(w242), .nr2(w242), .d(w248), .q(w1378) );
	dmg_dffr g351 (.clk(w476), .nr1(w242), .nr2(w242), .d(w1378), .q(w811) );
	dmg_dffr g352 (.clk(w476), .nr1(w242), .nr2(w242), .d(w811), .q(w477) );
	dmg_dffr g353 (.clk(w476), .nr1(w242), .nr2(w242), .d(w477), .q(w478) );
	dmg_dffr g354 (.clk(w809), .nr1(w1067), .nr2(w1067), .d(w1064), .q(w1267) );
	dmg_dffr g355 (.clk(w819), .nr1(w73), .nr2(w73), .d(w74), .q(w75), .nq(w74) );
	dmg_dffr g356 (.clk(w367), .nr1(w341), .nr2(w341), .d(w342), .q(w809) );
	dmg_dffr g357 (.clk(w162), .nr1(w152), .nr2(w152), .d(w303), .q(w151) );
	dmg_dffr g358 (.clk(w162), .nr1(w152), .nr2(w152), .d(w27), .q(w303) );
	dmg_dffr g359 (.clk(w162), .nr1(w918), .nr2(w918), .d(w919), .q(w27) );
	dmg_dffr g360 (.clk(w494), .nr1(w539), .nr2(w539), .d(w495), .q(w496), .nq(w495) );
	dmg_dffr g361 (.clk(w122), .nr1(w594), .nr2(w594), .d(w593), .q(w595) );
	dmg_dffr g362 (.clk(w654), .nr1(w656), .nr2(w656), .d(w657), .q(w658), .nq(w657) );
	dmg_dffr g363 (.clk(w1242), .nr1(w1320), .nr2(w1320), .d(w347), .q(w96) );
	dmg_dffr g364 (.clk(w122), .nr1(w1319), .nr2(w1319), .d(w1318), .q(w742) );
	dmg_dffr g365 (.clk(w282), .nr1(w1246), .nr2(w1246), .d(w404), .nq(w1245) );
	dmg_dffr g366 (.clk(w1207), .nr1(w40), .nr2(w40), .d(w41), .q(w925) );
	dmg_dffr g367 (.clk(w168), .nr1(w626), .nr2(w626), .d(w1292), .q(w914) );
	dmg_dffr g368 (.clk(w1092), .nr1(w818), .nr2(w818), .d(w149), .q(w220), .nq(w149) );
	dmg_dffr g369 (.clk(w279), .nr1(w818), .nr2(w818), .d(w1092), .q(w277), .nq(w1092) );
	dmg_dffr g370 (.clk(w1020), .nr1(w818), .nr2(w818), .d(w278), .q(w276), .nq(w278) );
	dmg_dffr g371 (.clk(w275), .nr1(w818), .nr2(w818), .d(w1020), .q(w1021), .nq(w1020) );
	dmg_dffr g372 (.clk(w1112), .nr1(w818), .nr2(w818), .d(w1058), .q(w1015), .nq(w1058) );
	dmg_dffr g373 (.clk(w1057), .nr1(w818), .nr2(w818), .d(w275), .q(w274), .nq(w275) );
	dmg_dffr g374 (.clk(w1391), .nr1(w818), .nr2(w818), .d(w1057), .q(w272), .nq(w1057) );
	dmg_dffr g375 (.clk(w1056), .nr1(w818), .nr2(w818), .d(w1391), .q(w841), .nq(w1391) );
	dmg_dffr g376 (.clk(w1055), .nr1(w818), .nr2(w818), .d(w1056), .q(w222), .nq(w1056) );
	dmg_dffr g377 (.clk(w283), .nr1(w1025), .nr2(w1025), .d(w1317), .nq(w1083) );
	dmg_dffr g378 (.clk(w1024), .nr1(w1025), .nr2(w1025), .d(w1084), .nq(w1084) );
	dmg_dffr g379 (.clk(w282), .nr1(w1134), .nr2(w1134), .d(w1023), .nq(w143) );
	dmg_dffr g380 (.clk(w282), .nr1(w307), .nr2(w307), .d(w308), .q(w292) );
	dmg_dffr g381 (.clk(w10), .nr1(w559), .nr2(w559), .d(w879), .q(w798) );
	dmg_dffr g382 (.clk(w1199), .nr1(w559), .nr2(w559), .d(w183), .q(w618) );
	dmg_dffr g383 (.clk(w709), .nr1(w19), .nr2(w19), .d(w16), .q(w86) );
	dmg_dffr g384 (.clk(w1166), .nr1(w696), .nr2(w696), .d(w86), .q(w85) );
	dmg_dffr g385 (.clk(w390), .nr1(w697), .nr2(w697), .d(w391), .q(w392) );
	dmg_dffr g386 (.clk(w388), .nr1(w697), .nr2(w697), .d(w659), .q(w391) );
	dmg_cnt g387 (.d(w16), .load(w708), .nq(w1167), .clk(w1160) );
	dmg_cnt g388 (.q(w1022), .d(w940), .load(w1028), .clk(w280) );
	dmg_cnt g389 (.q(w1081), .d(w1080), .load(w1028), .clk(w1022) );
	dmg_cnt g390 (.q(w288), .d(w941), .load(w1316), .clk(w290) );
	dmg_cnt g391 (.q(w290), .d(w309), .load(w1316), .clk(w289) );
	dmg_cnt g392 (.q(w289), .d(w1076), .load(w1316), .clk(w287) );
	dmg_cnt g393 (.d(w229), .load(w321), .nq(w286), .clk(w82) );
	dmg_cnt g394 (.q(w1190), .d(w305), .load(w913), .nq(w825), .clk(w153) );
	dmg_cnt g395 (.q(w996), .d(w1119), .load(w968), .clk(w1034) );
	dmg_cnt g396 (.q(w1034), .d(w967), .load(w968), .clk(w950) );
	dmg_cnt g397 (.q(w954), .d(w331), .load(w952), .clk(w1329) );
	dmg_cnt g398 (.d(w229), .load(w952), .nq(w963), .clk(w953) );
	dmg_cnt g399 (.q(w1263), .d(w29), .load(w1264), .clk(w1302) );
	dmg_cnt g400 (.q(w1171), .d(w331), .load(w571), .clk(w1170) );
	dmg_cnt g401 (.q(w759), .d(w180), .load(w571), .clk(w1171) );
	dmg_cnt g402 (.d(w229), .load(w571), .nq(w758), .clk(w759) );
	dmg_cnt g403 (.d(w750), .load(w646), .nq(w1212), .clk(w1238) );
	dmg_cnt g404 (.q(w1238), .d(w1239), .load(w646), .nq(w1240), .clk(w653) );
	dmg_cnt g405 (.q(w1170), .d(w183), .load(w571), .clk(w1174) );
	dmg_cnt g406 (.d(w16), .load(w1264), .nq(w1265), .clk(w1263) );
	dmg_cnt g407 (.d(w997), .load(w160), .nq(w912), .clk(w159) );
	dmg_cnt g408 (.q(w1115), .d(w297), .load(w913), .nq(w911), .clk(w910) );
	dmg_cnt g409 (.q(w153), .d(w931), .load(w913), .nq(w1005), .clk(w1115) );
	dmg_cnt g410 (.d(w16), .load(w319), .nq(w819), .clk(w852) );
	dmg_cnt g411 (.q(w330), .d(w860), .load(w845), .nq(w326), .clk(w325) );
	dmg_cnt g412 (.d(w229), .load(w916), .nq(w1278), .clk(w540) );
	dmg_cnt g413 (.q(w540), .d(w180), .load(w916), .clk(w1373) );
	dmg_cnt g414 (.q(w1279), .d(w183), .load(w916), .clk(w1280) );
	dmg_cnt g415 (.q(w536), .d(w29), .load(w170), .clk(w1277) );
	dmg_cnt g416 (.d(w1357), .load(w550), .nq(w525), .clk(w1338) );
	dmg_cnt g417 (.q(w1336), .d(w1337), .load(w550), .nq(w1321), .clk(w1322) );
	dmg_cnt g418 (.q(w1338), .d(w549), .load(w550), .nq(w739), .clk(w1336) );
	dmg_cnt g419 (.q(w602), .d(w736), .load(w735), .nq(w1258), .clk(w173) );
	dmg_cnt g420 (.q(w605), .d(w633), .load(w365), .clk(w732) );
	dmg_cnt g421 (.q(w732), .d(w364), .load(w365), .clk(w676) );
	dmg_cnt g422 (.q(w676), .d(w729), .load(w365), .clk(w727) );
	dmg_cnt g423 (.q(w1234), .d(w1228), .load(w371), .clk(w1222) );
	dmg_cnt g424 (.q(w534), .d(w254), .load(w160), .nq(w1128), .clk(w255) );
	dmg_cnt g425 (.q(w257), .d(w567), .load(w845), .nq(w569), .clk(w568) );
	dmg_cnt g426 (.q(w1369), .d(w138), .load(w137), .clk(w1014) );
	dmg_cnt g427 (.q(w333), .d(w332), .load(w137), .clk(w1369) );
	dmg_cnt g428 (.q(w1368), .d(w1272), .load(w137), .clk(w333) );
	dmg_cnt g429 (.d(w566), .load(w845), .nq(w256), .clk(w257) );
	dmg_cnt g430 (.q(w373), .d(w1283), .load(w371), .clk(w1234) );
	dmg_cnt g431 (.q(w372), .d(w374), .load(w371), .clk(w373) );
	dmg_cnt g432 (.q(w446), .d(w199), .load(w198), .nq(w178), .clk(w179) );
	dmg_cnt g433 (.q(w179), .d(w448), .load(w198), .nq(w447), .clk(w445) );
	dmg_cnt g434 (.d(w731), .load(w198), .nq(w462), .clk(w446) );
	dmg_cnt g435 (.q(w445), .d(w449), .load(w198), .nq(w634), .clk(w604) );
	dmg_cnt g436 (.q(w635), .d(w464), .load(w196), .nq(w459), .clk(w460) );
	dmg_cnt g437 (.q(w460), .d(w195), .load(w196), .nq(w636), .clk(w463) );
	dmg_cnt g438 (.q(w463), .d(w193), .load(w196), .nq(w192), .clk(w461) );
	dmg_cnt g439 (.d(w375), .load(w196), .nq(w186), .clk(w635) );
	dmg_cnt g440 (.q(w1388), .d(w734), .load(w735), .nq(w184), .clk(w185) );
	dmg_cnt g441 (.q(w173), .d(w1286), .load(w735), .nq(w1287), .clk(w1388) );
	dmg_cnt g442 (.q(w1382), .d(w455), .load(w456), .nq(w608), .clk(w607) );
	dmg_cnt g443 (.q(w607), .d(w606), .load(w456), .nq(w1351), .clk(w1352) );
	dmg_cnt g444 (.q(w1352), .d(w457), .load(w456), .nq(w908), .clk(w552) );
	dmg_cnt g445 (.q(w440), .d(w438), .load(w27), .nq(w441), .clk(w442) );
	dmg_cnt g446 (.q(w471), .d(w530), .load(w27), .clk(w847) );
	dmg_cnt g447 (.q(w541), .d(w848), .load(w27), .nq(w533), .clk(w157) );
	dmg_cnt g448 (.q(w158), .d(w874), .load(w160), .nq(w535), .clk(w534) );
	dmg_cnt g449 (.q(w156), .d(w214), .load(w27), .nq(w532), .clk(w531) );
	dmg_cnt g450 (.q(w568), .d(w789), .load(w845), .nq(w329), .clk(w330) );
	dmg_cnt g451 (.q(w1061), .d(w480), .load(w340), .nq(w1268), .clk(w1063) );
	dmg_cnt g452 (.q(w834), .d(w481), .load(w340), .clk(w1062) );
	dmg_cnt g453 (.q(w129), .d(w339), .load(w340), .nq(w1060), .clk(w835) );
	dmg_cnt g454 (.q(w133), .d(w1269), .load(w340), .nq(w980), .clk(w617) );
	dmg_cnt g455 (.q(w852), .d(w29), .load(w319), .clk(w285) );
	dmg_cnt g456 (.q(w81), .d(w331), .load(w321), .clk(w80) );
	dmg_cnt g457 (.q(w159), .d(w764), .load(w160), .nq(w1191), .clk(w158) );
	dmg_cnt g458 (.q(w1373), .d(w331), .load(w916), .clk(w1279) );
	dmg_cnt g459 (.d(w187), .load(w170), .nq(w494), .clk(w171) );
	dmg_cnt g460 (.q(w171), .d(w55), .load(w170), .clk(w1393) );
	dmg_cnt g461 (.q(w1393), .d(w16), .load(w170), .clk(w536) );
	dmg_cnt g462 (.q(w353), .d(w352), .load(w347), .nq(w899), .clk(w900) );
	dmg_cnt g463 (.q(w91), .d(w351), .load(w347), .nq(w897), .clk(w898) );
	dmg_cnt g464 (.q(w355), .d(w348), .load(w347), .nq(w356), .clk(w357) );
	dmg_cnt g465 (.q(w1209), .d(w361), .load(w347), .clk(w362) );
	dmg_cnt g466 (.q(w1322), .d(w1289), .load(w550), .nq(w1323), .clk(w1213) );
	dmg_cnt g467 (.q(w741), .d(w748), .load(w646), .nq(w747), .clk(w101) );
	dmg_cnt g468 (.q(w653), .d(w652), .load(w646), .nq(w740), .clk(w741) );
	dmg_cnt g469 (.q(w995), .d(w994), .load(w968), .clk(w996) );
	dmg_cnt g470 (.q(w82), .d(w180), .load(w321), .clk(w81) );
	dmg_cnt g471 (.q(w80), .d(w183), .load(w321), .clk(w79) );
	dmg_cnt g472 (.q(w1082), .d(w1090), .load(w1028), .clk(w1081) );
	dmg_cnt g473 (.q(w1329), .d(w183), .load(w952), .clk(w1294) );
	dmg_cnt g474 (.q(w953), .d(w180), .load(w952), .clk(w954) );
	dmg_cnt g475 (.q(w1160), .d(w29), .load(w708), .clk(w1333) );
	dmg_latchr_comp g476 (.n_ena(w230), .d(w29), .ena(w142), .nres(w942), .nq(w1076) );
	dmg_latchr_comp g477 (.n_ena(w230), .d(w229), .ena(w142), .nres(w942), .nq(w1079) );
	dmg_latchr_comp g478 (.n_ena(w230), .d(w180), .ena(w142), .nres(w942), .nq(w1090) );
	dmg_latchr_comp g479 (.n_ena(w230), .d(w331), .ena(w142), .nres(w942), .nq(w1080) );
	dmg_latchr_comp g480 (.n_ena(w1104), .d(w183), .ena(w988), .nres(w19), .q(w18), .nq(w1154) );
	dmg_latchr_comp g481 (.n_ena(w1104), .d(w229), .ena(w988), .nres(w19), .q(w17), .nq(w813) );
	dmg_latchr_comp g482 (.n_ena(w1103), .d(w183), .ena(w228), .nres(w19), .nq(w227) );
	dmg_latchr_comp g483 (.n_ena(w1103), .d(w229), .ena(w228), .nres(w19), .q(w815), .nq(w814) );
	dmg_latchr_comp g484 (.n_ena(w1103), .d(w180), .ena(w228), .nres(w19), .nq(w1153) );
	dmg_latchr_comp g485 (.n_ena(w1074), .d(w55), .ena(w1075), .nres(w19), .nq(w224) );
	dmg_latchr_comp g486 (.n_ena(w69), .d(w55), .ena(w1107), .nres(w1106), .q(w76), .nq(w77) );
	dmg_latchr_comp g487 (.n_ena(w625), .d(w55), .ena(w624), .nres(w626), .q(w485), .nq(w484) );
	dmg_latchr_comp g488 (.n_ena(w753), .d(w403), .ena(w379), .nres(w519), .nq(w751) );
	dmg_latchr_comp g489 (.n_ena(w753), .d(w1157), .ena(w379), .nres(w519), .nq(w752) );
	dmg_latchr_comp g490 (.n_ena(w515), .d(w514), .ena(w379), .nres(w519), .nq(w522) );
	dmg_latchr_comp g491 (.n_ena(w515), .d(w380), .ena(w379), .nres(w519), .nq(w1247) );
	dmg_latchr_comp g492 (.n_ena(w1172), .d(w187), .ena(w1150), .nres(w1384), .q(w1318) );
	dmg_latchr_comp g493 (.n_ena(w510), .d(w55), .ena(w511), .nres(w509), .q(w508), .nq(w506) );
	dmg_latchr_comp g494 (.n_ena(w1180), .d(w331), .ena(w1179), .nres(w338), .q(w1118), .nq(w1119) );
	dmg_latchr_comp g495 (.n_ena(w1180), .d(w180), .ena(w1179), .nres(w338), .q(w1182), .nq(w994) );
	dmg_latchr_comp g496 (.n_ena(w1180), .d(w183), .ena(w1179), .nres(w338), .q(w1117), .nq(w967) );
	dmg_latchr_comp g497 (.n_ena(w337), .d(w55), .ena(w810), .nres(w338), .q(w480), .nq(w54) );
	dmg_latchr_comp g498 (.n_ena(w337), .d(w16), .ena(w810), .nres(w338), .q(w339), .nq(w1370) );
	dmg_latchr_comp g499 (.n_ena(w337), .d(w187), .ena(w810), .nres(w338), .q(w481), .nq(w482) );
	dmg_latchr_comp g500 (.n_ena(w337), .d(w229), .ena(w810), .nres(w338), .q(w134), .nq(w616) );
	dmg_latchr_comp g501 (.n_ena(w337), .d(w29), .ena(w810), .nres(w338), .q(w1269), .nq(w1270) );
	dmg_latchr_comp g502 (.n_ena(w974), .d(w55), .ena(w975), .nres(w818), .q(w1016), .nq(w1111) );
	dmg_latchr_comp g503 (.n_ena(w974), .d(w187), .ena(w975), .nres(w818), .q(w973), .nq(w475) );
	dmg_latchr_comp g504 (.n_ena(w1193), .d(w187), .ena(w1194), .nres(w1192), .q(w409), .nq(w408) );
	dmg_latchr_comp g505 (.n_ena(w722), .d(w16), .ena(w1211), .nres(w363), .q(w351), .nq(w350) );
	dmg_latchr_comp g506 (.n_ena(w722), .d(w55), .ena(w1211), .nres(w363), .q(w348), .nq(w349) );
	dmg_latchr_comp g507 (.n_ena(w722), .d(w29), .ena(w1211), .nres(w363), .q(w352), .nq(w557) );
	dmg_latchr_comp g508 (.n_ena(w722), .d(w187), .ena(w1211), .nres(w363), .q(w361), .nq(w360) );
	dmg_latchr_comp g509 (.n_ena(w548), .d(w187), .ena(w1251), .nres(w749), .q(w1357) );
	dmg_latchr_comp g510 (.n_ena(w548), .d(w55), .ena(w1251), .nres(w749), .q(w549) );
	dmg_latchr_comp g511 (.n_ena(w548), .d(w16), .ena(w1251), .nres(w749), .q(w1337) );
	dmg_latchr_comp g512 (.n_ena(w553), .d(w187), .ena(w554), .nres(w592), .q(w593) );
	dmg_latchr_comp g513 (.n_ena(w182), .d(w331), .ena(w181), .nres(w197), .q(w1286) );
	dmg_latchr_comp g514 (.n_ena(w182), .d(w183), .ena(w181), .nres(w197), .q(w734) );
	dmg_latchr_comp g515 (.n_ena(w182), .d(w180), .ena(w181), .nres(w197), .q(w736) );
	dmg_latchr_comp g516 (.n_ena(w450), .d(w183), .ena(w451), .nres(w458), .q(w457) );
	dmg_latchr_comp g517 (.n_ena(w450), .d(w180), .ena(w451), .nres(w458), .q(w455) );
	dmg_latchr_comp g518 (.n_ena(w450), .d(w331), .ena(w451), .nres(w458), .q(w606) );
	dmg_latchr_comp g519 (.n_ena(w201), .d(w331), .ena(w200), .nres(w194), .q(w448) );
	dmg_latchr_comp g520 (.n_ena(w201), .d(w29), .ena(w200), .nres(w194), .q(w193) );
	dmg_latchr_comp g521 (.n_ena(w201), .d(w229), .ena(w200), .nres(w194), .q(w731) );
	dmg_latchr_comp g522 (.n_ena(w201), .d(w180), .ena(w200), .nres(w194), .q(w199) );
	dmg_latchr_comp g523 (.n_ena(w202), .d(w16), .ena(w203), .nres(w194), .q(w195) );
	dmg_latchr_comp g524 (.n_ena(w1227), .d(w183), .ena(w724), .nres(w430), .q(w1285), .nq(w1228) );
	dmg_latchr_comp g525 (.n_ena(w1227), .d(w180), .ena(w724), .nres(w430), .q(w429), .nq(w374) );
	dmg_latchr_comp g526 (.n_ena(w1227), .d(w331), .ena(w724), .nres(w430), .q(w1284), .nq(w1283) );
	dmg_latchr_comp g527 (.n_ena(w851), .d(w16), .ena(w1282), .nres(w430), .q(w214), .nq(w213) );
	dmg_latchr_comp g528 (.n_ena(w851), .d(w29), .ena(w1282), .nres(w430), .q(w438), .nq(w850) );
	dmg_latchr_comp g529 (.n_ena(w851), .d(w55), .ena(w1282), .nres(w430), .q(w848), .nq(w849) );
	dmg_latchr_comp g530 (.n_ena(w851), .d(w229), .ena(w1282), .nres(w430), .q(w439), .nq(w433) );
	dmg_latchr_comp g531 (.n_ena(w851), .d(w187), .ena(w1282), .nres(w430), .q(w530), .nq(w431) );
	dmg_latchr_comp g532 (.n_ena(w1377), .d(w331), .ena(w1271), .nres(w139), .nq(w332) );
	dmg_latchr_comp g533 (.n_ena(w1377), .d(w180), .ena(w1271), .nres(w139), .nq(w1272) );
	dmg_latchr_comp g534 (.n_ena(w1377), .d(w183), .ena(w1271), .nres(w139), .nq(w138) );
	dmg_latchr_comp g535 (.n_ena(w334), .d(w229), .ena(w335), .nres(w52), .q(w783), .nq(w782) );
	dmg_latchr_comp g536 (.n_ena(w202), .d(w55), .ena(w203), .nres(w194), .q(w464) );
	dmg_latchr_comp g537 (.n_ena(w202), .d(w187), .ena(w203), .nres(w194), .q(w375) );
	dmg_latchr_comp g538 (.n_ena(w201), .d(w183), .ena(w200), .nres(w194), .q(w449) );
	dmg_latchr_comp g539 (.n_ena(w1356), .d(w16), .ena(w1355), .nres(w1354), .q(w591), .nq(w588) );
	dmg_latchr_comp g540 (.n_ena(w1356), .d(w55), .ena(w1355), .nres(w1354), .q(w589), .nq(w590) );
	dmg_latchr_comp g541 (.n_ena(w675), .d(w331), .ena(w674), .nres(w363), .q(w1257), .nq(w364) );
	dmg_latchr_comp g542 (.n_ena(w675), .d(w180), .ena(w674), .nres(w363), .q(w1256), .nq(w633) );
	dmg_latchr_comp g543 (.n_ena(w675), .d(w183), .ena(w674), .nres(w363), .q(w728), .nq(w729) );
	dmg_latchr_comp g544 (.n_ena(w537), .d(w55), .ena(w538), .nres(w1217), .q(w497), .nq(w498) );
	dmg_latchr_comp g545 (.n_ena(w821), .d(w187), .ena(w1358), .nres(w261), .q(w260) );
	dmg_latchr_comp g546 (.n_ena(w974), .d(w29), .ena(w975), .nres(w818), .q(w982), .nq(w971) );
	dmg_latchr_comp g547 (.n_ena(w974), .d(w16), .ena(w975), .nres(w818), .q(w983), .nq(w972) );
	dmg_latchr_comp g548 (.n_ena(w722), .d(w229), .ena(w1211), .nres(w363), .q(w502), .nq(w358) );
	dmg_latchr_comp g549 (.n_ena(w1250), .d(w1252), .ena(w638), .nres(w19), .q(w1029), .nq(w1210) );
	dmg_latchr_comp g550 (.n_ena(w651), .d(w29), .ena(w650), .nres(w749), .q(w1289) );
	dmg_latchr_comp g551 (.n_ena(w651), .d(w229), .ena(w650), .nres(w749), .q(w750) );
	dmg_latchr_comp g552 (.n_ena(w651), .d(w180), .ena(w650), .nres(w749), .q(w1239) );
	dmg_latchr_comp g553 (.n_ena(w651), .d(w331), .ena(w650), .nres(w749), .q(w652) );
	dmg_latchr_comp g554 (.n_ena(w651), .d(w183), .ena(w650), .nres(w749), .q(w748) );
	dmg_latchr_comp g555 (.n_ena(w625), .d(w187), .ena(w624), .nres(w626), .q(w629), .nq(w630) );
	dmg_latchr_comp g556 (.n_ena(w1006), .d(w187), .ena(w1007), .nres(w921), .q(w922) );
	dmg_latchr_comp g557 (.n_ena(w1103), .d(w331), .ena(w228), .nres(w19), .nq(w376) );
	dmg_latchr_comp g558 (.n_ena(w1104), .d(w331), .ena(w988), .nres(w19), .q(w1108), .nq(w1105) );
	dmg_latchr_comp g559 (.n_ena(w1104), .d(w180), .ena(w988), .nres(w19), .q(w816), .nq(w817) );
	dmg_latchr_comp g560 (.n_ena(w1074), .d(w16), .ena(w1075), .nres(w19), .nq(w1151) );
	dmg_latchr_comp g561 (.n_ena(w1074), .d(w187), .ena(w1075), .nres(w19), .q(w1109), .nq(w1110) );
	dmg_latchr_comp g562 (.n_ena(w1074), .d(w29), .ena(w1075), .nres(w19), .nq(w226) );
	dmg_latchr_comp g563 (.n_ena(w191), .d(w16), .ena(w190), .nres(w19), .q(w1072), .nq(w1073) );
	dmg_latchr_comp g564 (.n_ena(w191), .d(w29), .ena(w190), .nres(w19), .q(w1094), .nq(w1093) );
	dmg_latchr_comp g565 (.n_ena(w191), .d(w55), .ena(w190), .nres(w19), .q(w1047), .nq(w840) );
	dmg_latchr_comp g566 (.n_ena(w191), .d(w187), .ena(w190), .nres(w19), .q(w1048), .nq(w1049) );
	dmg_latchr_comp g567 (.n_ena(w230), .d(w16), .ena(w142), .nres(w942), .nq(w309) );
	dmg_latchr_comp g568 (.n_ena(w230), .d(w183), .ena(w142), .nres(w942), .nq(w940) );
	dmg_latchr_comp g569 (.n_ena(w230), .d(w55), .ena(w142), .nres(w942), .nq(w941) );
	dmg_latchr_comp g570 (.n_ena(w944), .d(w55), .ena(w945), .nres(w946), .q(w23), .nq(w1100) );
	dmg_latchr_comp g571 (.n_ena(w663), .d(w55), .ena(w1122), .nres(w40), .q(w34), .nq(w35) );
	dmg_latchr_comp g572 (.n_ena(w663), .d(w187), .ena(w1122), .nres(w40), .q(w37), .nq(w36) );
	dmg_latchr_comp g573 (.n_ena(w378), .d(w583), .ena(w379), .nres(w519), .nq(w585) );
	dmg_latchr_comp g574 (.n_ena(w378), .d(w584), .ena(w379), .nres(w519), .nq(w520) );
	dmg_latchr_comp g575 (.n_ena(w516), .d(w573), .ena(w379), .nres(w519), .nq(w518) );
	dmg_latchr_comp g576 (.n_ena(w516), .d(w1162), .ena(w379), .nres(w519), .nq(w517) );
	dmg_nor g577 (.a(w90), .b(w3), .x(w2) );
	dmg_not2 g578 (.a(w104), .x(w206) );
	dmg_not2 g579 (.a(w103), .x(w62) );
	dmg_not2 g580 (.a(w110), .x(w208) );
	dmg_nor g581 (.a(w755), .b(w70), .x(w959) );
	dmg_not2 g582 (.a(w12), .x(w13) );
	dmg_nor g583 (.a(w90), .b(w13), .x(w14) );
	dmg_nor g584 (.a(w546), .b(w70), .x(w1308) );
	dmg_nor g585 (.a(w70), .b(w1312), .x(w1315) );
	dmg_nor g586 (.a(w70), .b(w1045), .x(w1327) );
	dmg_nor g587 (.a(w70), .b(w1350), .x(w1311) );
	dmg_nor g588 (.a(w70), .b(w292), .x(w1134) );
	dmg_nor g589 (.a(w44), .b(w312), .x(w311) );
	dmg_nor g590 (.a(w1248), .b(w887), .x(w886) );
	dmg_nor g591 (.a(w1036), .b(w887), .x(w1035) );
	dmg_nor g592 (.a(w484), .b(w629), .x(w1301) );
	dmg_nor g593 (.a(w485), .b(w629), .x(w628) );
	dmg_nor g594 (.a(w485), .b(w630), .x(w486) );
	dmg_nor g595 (.a(w484), .b(w630), .x(w1300) );
	dmg_nor g596 (.a(w1041), .b(w887), .x(w824) );
	dmg_nor g597 (.a(w990), .b(w887), .x(w823) );
	dmg_nor g598 (.a(w453), .b(w61), .x(w60) );
	dmg_nor g599 (.a(w90), .b(w1123), .x(w89) );
	dmg_nor g600 (.a(w453), .b(w205), .x(w204) );
	dmg_nor g601 (.a(w90), .b(w1331), .x(w621) );
	dmg_not2 g602 (.a(w1245), .x(w397) );
	dmg_nor g603 (.a(w90), .b(w1237), .x(w1244) );
	dmg_nor g604 (.a(w1242), .b(w99), .x(w100) );
	dmg_nor g605 (.a(w346), .b(w658), .x(w108) );
	dmg_nor g606 (.a(w453), .b(w641), .x(w401) );
	dmg_nor g607 (.a(w453), .b(w402), .x(w210) );
	dmg_nor g608 (.a(w1324), .b(w70), .x(w1214) );
	dmg_nor g609 (.a(w762), .b(w70), .x(w1325) );
	dmg_nor g610 (.a(w761), .b(w70), .x(w414) );
	dmg_nor g611 (.a(w70), .b(w303), .x(w918) );
	dmg_nor g612 (.a(w168), .b(w27), .x(w161) );
	dmg_nor g613 (.a(w70), .b(w1116), .x(w1185) );
	dmg_nor g614 (.a(w70), .b(w869), .x(w870) );
	dmg_nor g615 (.a(w292), .b(w151), .x(w150) );
	dmg_nor g616 (.a(w70), .b(w144), .x(w145) );
	dmg_nor g617 (.a(w340), .b(w809), .x(w969) );
	dmg_nor g618 (.a(w146), .b(w162), .x(w147) );
	dmg_nor g619 (.a(w340), .b(w70), .x(w1067) );
	dmg_nor g620 (.a(w70), .b(w340), .x(w479) );
	dmg_nor g621 (.a(w340), .b(w271), .x(w136) );
	dmg_nor g622 (.a(w70), .b(w120), .x(w261) );
	dmg_nor g623 (.a(w976), .b(w70), .x(w1374) );
	dmg_nor g624 (.a(w528), .b(w70), .x(w472) );
	dmg_nor g625 (.a(w328), .b(w70), .x(w215) );
	dmg_nor g626 (.a(w720), .b(w453), .x(w454) );
	dmg_nor g627 (.a(w905), .b(w610), .x(w719) );
	dmg_nor g628 (.a(w906), .b(w175), .x(w176) );
	dmg_nor g629 (.a(w589), .b(w588), .x(w524) );
	dmg_nor g630 (.a(w590), .b(w591), .x(w649) );
	dmg_nor g631 (.a(w590), .b(w588), .x(w587) );
	dmg_nor g632 (.a(w70), .b(w250), .x(w269) );
	dmg_nor g633 (.a(w27), .b(w70), .x(w425) );
	dmg_nor g634 (.a(w70), .b(w240), .x(w239) );
	dmg_nor g635 (.a(w292), .b(w27), .x(w233) );
	dmg_nor g636 (.a(w70), .b(w238), .x(w216) );
	dmg_nor g637 (.a(w619), .b(w563), .x(w876) );
	dmg_nor g638 (.a(w367), .b(w368), .x(w1380) );
	dmg_nor g639 (.a(w560), .b(w563), .x(w561) );
	dmg_nor g640 (.a(w27), .b(w369), .x(w370) );
	dmg_nor g641 (.a(w1274), .b(w70), .x(w418) );
	dmg_nor g642 (.a(w1127), .b(w70), .x(w936) );
	dmg_nor g643 (.a(w846), .b(w563), .x(w564) );
	dmg_nor g644 (.a(w1381), .b(w563), .x(w938) );
	dmg_nor g645 (.a(w90), .b(w128), .x(w127) );
	dmg_nor g646 (.a(w1230), .b(w1126), .x(w1273) );
	dmg_nor g647 (.a(w1231), .b(w803), .x(w802) );
	dmg_nor g648 (.a(w686), .b(w685), .x(w603) );
	dmg_nor g649 (.a(w659), .b(w346), .x(w345) );
	dmg_nor g650 (.a(w347), .b(w70), .x(w95) );
	dmg_nor g651 (.a(w347), .b(w679), .x(w366) );
	dmg_nor g652 (.a(w367), .b(w680), .x(w672) );
	dmg_nor g653 (.a(w367), .b(w808), .x(w856) );
	dmg_nor g654 (.a(w70), .b(w1379), .x(w864) );
	dmg_nor g655 (.a(w70), .b(w791), .x(w785) );
	dmg_nor g656 (.a(w836), .b(w70), .x(w1361) );
	dmg_nor g657 (.a(w44), .b(w473), .x(w53) );
	dmg_nor g658 (.a(w70), .b(w71), .x(w853) );
	dmg_nor g659 (.a(w162), .b(w323), .x(w324) );
	dmg_nor g660 (.a(w529), .b(w70), .x(w322) );
	dmg_nor g661 (.a(w639), .b(w453), .x(w452) );
	dmg_nor g662 (.a(w408), .b(w70), .x(w344) );
	dmg_nor g663 (.a(w70), .b(w595), .x(w592) );
	dmg_nor g664 (.a(w70), .b(w599), .x(w598) );
	dmg_nor g665 (.a(w70), .b(w96), .x(w744) );
	dmg_nor g666 (.a(w70), .b(w742), .x(w1384) );
	dmg_nor g667 (.a(w453), .b(w1173), .x(w904) );
	dmg_nor g668 (.a(w453), .b(w1149), .x(w504) );
	dmg_nor g669 (.a(w503), .b(w453), .x(w501) );
	dmg_nor g670 (.a(w453), .b(w903), .x(w902) );
	dmg_nor g671 (.a(w1207), .b(w347), .x(w551) );
	dmg_nor g672 (.a(w35), .b(w37), .x(w1291) );
	dmg_nor g673 (.a(w34), .b(w37), .x(w33) );
	dmg_nor g674 (.a(w35), .b(w36), .x(w894) );
	dmg_nor g675 (.a(w34), .b(w36), .x(w888) );
	dmg_nor g676 (.a(w642), .b(w453), .x(w1297) );
	dmg_nor g677 (.a(w453), .b(w314), .x(w313) );
	dmg_nor g678 (.a(w453), .b(w64), .x(w65) );
	dmg_nor g679 (.a(w453), .b(w991), .x(w943) );
	dmg_nor g680 (.a(w962), .b(w887), .x(w1218) );
	dmg_nor g681 (.a(w66), .b(w67), .x(w343) );
	dmg_nor g682 (.a(w70), .b(w920), .x(w921) );
	dmg_nor g683 (.a(w292), .b(w27), .x(w291) );
	dmg_nor g684 (.a(w27), .b(w292), .x(w1027) );
	dmg_nor g685 (.a(w1026), .b(w147), .x(w148) );
	dmg_nor g686 (.a(w1133), .b(w70), .x(w307) );
	dmg_nor g687 (.a(w231), .b(w1086), .x(w1087) );
	dmg_nor g688 (.a(w70), .b(w1314), .x(w999) );
	dmg_nor g689 (.a(w1346), .b(w70), .x(w1183) );
	dmg_nor g690 (.a(w1349), .b(w70), .x(w296) );
	dmg_nor g691 (.a(w44), .b(w1097), .x(w1096) );
	dmg_nor g692 (.a(w1201), .b(w1198), .x(w695) );
	dmg_nor g693 (.a(w1198), .b(w665), .x(w664) );
	dmg_nor g694 (.a(w90), .b(w694), .x(w622) );
	dmg_nor g695 (.a(w90), .b(w693), .x(w1040) );
	dmg_nor g696 (.a(w90), .b(w662), .x(w661) );
	dmg_nor g697 (.a(w393), .b(w394), .x(w395) );
	dmg_not3 g698 (.a(w1164), .x(w1163) );
	dmg_not3 g699 (.a(w1332), .x(w705) );
	dmg_not3 g700 (.a(w574), .x(w575) );
	dmg_not3 g701 (.a(w1084), .x(w1042) );
	dmg_not3 g702 (.a(w1079), .x(w231) );
	dmg_not3 g703 (.a(w1024), .x(w1188) );
	dmg_not3 g704 (.a(w1206), .x(w582) );
	dmg_not3 g705 (.a(w218), .x(w217) );
	dmg_not3 g706 (.a(w148), .x(w219) );
	dmg_not3 g707 (.a(w774), .x(w19) );
	dmg_not3 g708 (.a(w857), .x(w367) );
	dmg_not3 g709 (.a(w284), .x(w263) );
	dmg_not3 g710 (.a(w1307), .x(w1043) );
	dmg_not3 g711 (.a(w1304), .x(w1008) );
	dmg_not3 g712 (.a(w1295), .x(w957) );
	dmg_not2 g713 (.a(w14), .x(w15) );
	dmg_not2 g714 (.a(w142), .x(w230) );
	dmg_not2 g715 (.a(w311), .x(w310) );
	dmg_not2 g716 (.a(w190), .x(w191) );
	dmg_not2 g717 (.a(w1096), .x(w225) );
	dmg_not2 g718 (.a(w988), .x(w1104) );
	dmg_not2 g719 (.a(w228), .x(w1103) );
	dmg_not2 g720 (.a(w650), .x(w651) );
	dmg_not2 g721 (.a(w1211), .x(w722) );
	dmg_not2 g722 (.a(w343), .x(w28) );
	dmg_not2 g723 (.a(w975), .x(w974) );
	dmg_not2 g724 (.a(w53), .x(w812) );
	dmg_not2 g725 (.a(w1181), .x(w242) );
	dmg_not2 g726 (.a(w437), .x(w298) );
	dmg_not2 g727 (.a(w1282), .x(w851) );
	dmg_not2 g728 (.a(w200), .x(w201) );
	dmg_not2 g729 (.a(w176), .x(w177) );
	dmg_not2 g730 (.a(w559), .x(w1130) );
	dmg_not2 g731 (.a(w1271), .x(w1377) );
	dmg_not2 g732 (.a(w810), .x(w337) );
	dmg_not2 g733 (.a(w719), .x(w526) );
	dmg_not2 g734 (.a(w208), .x(w640) );
	dmg_not2 g735 (.a(w206), .x(w315) );
	dmg_not2 g736 (.a(w62), .x(w63) );
	dmg_not2 g737 (.a(w209), .x(w207) );
	dmg_not2 g738 (.a(w667), .x(w209) );
	dmg_not2 g739 (.a(w295), .x(w162) );
	dmg_not2 g740 (.a(w70), .x(w818) );
	dmg_not2 g741 (.a(w698), .x(w379) );
	dmg_not2 g742 (.a(w580), .x(w581) );
	dmg_not2 g743 (.a(w664), .x(w453) );
	dmg_not2 g744 (.a(w189), .x(w988) );
	dmg_not2 g745 (.a(w189), .x(w190) );
	dmg_not2 g746 (.a(w1083), .x(w284) );
	dmg_not2 g747 (.a(w1102), .x(w228) );
	dmg_not2 g748 (.a(w1102), .x(w1075) );
	dmg_not2 g749 (.a(w1075), .x(w1074) );
	dmg_nand g750 (.a(w188), .b(w204), .x(w1158) );
	dmg_nand g751 (.a(w180), .b(w294), .x(w1309) );
	dmg_nand g752 (.a(w1331), .b(w125), .x(w701) );
	dmg_nand g753 (.a(w1237), .b(w125), .x(w1243) );
	dmg_nand g754 (.a(w188), .b(w501), .x(w553) );
	dmg_nand g755 (.a(w1120), .b(w611), .x(w175) );
	dmg_nand g756 (.a(w55), .b(w30), .x(w558) );
	dmg_nand g757 (.a(w187), .b(w30), .x(w172) );
	dmg_nand g758 (.a(w631), .b(w504), .x(w510) );
	dmg_nand g759 (.a(w764), .b(w236), .x(w302) );
	dmg_nand g760 (.a(w874), .b(w236), .x(w264) );
	dmg_nand g761 (.a(w229), .b(w30), .x(w884) );
	dmg_nand g762 (.a(w183), .b(w30), .x(w1114) );
	dmg_nand g763 (.a(w180), .b(w30), .x(w788) );
	dmg_nand g764 (.a(w331), .b(w30), .x(w259) );
	dmg_nand g765 (.a(w501), .b(w500), .x(w499) );
	dmg_nand g766 (.a(w1335), .b(w637), .x(w1254) );
	dmg_nand g767 (.a(w336), .b(w42), .x(w909) );
	dmg_nand g768 (.a(w637), .b(w1392), .x(w47) );
	dmg_nand g769 (.a(w566), .b(w236), .x(w796) );
	dmg_nand g770 (.a(w254), .b(w236), .x(w253) );
	dmg_nand g771 (.a(w619), .b(w618), .x(w435) );
	dmg_nand g772 (.a(w560), .b(w618), .x(w877) );
	dmg_nand g773 (.a(w29), .b(w30), .x(w417) );
	dmg_nand g774 (.a(w16), .b(w30), .x(w1326) );
	dmg_nand g775 (.a(w846), .b(w618), .x(w937) );
	dmg_nand g776 (.a(w1381), .b(w618), .x(w939) );
	dmg_nand g777 (.a(w128), .b(w125), .x(w126) );
	dmg_nand g778 (.a(w1126), .b(w881), .x(w882) );
	dmg_nand g779 (.a(w803), .b(w618), .x(w804) );
	dmg_nand g780 (.a(w454), .b(w730), .x(w907) );
	dmg_nand g781 (.a(w637), .b(w188), .x(w1255) );
	dmg_nand g782 (.a(w504), .b(w1221), .x(w505) );
	dmg_nand g783 (.a(w567), .b(w234), .x(w1371) );
	dmg_nand g784 (.a(w789), .b(w234), .x(w235) );
	dmg_nand g785 (.a(w860), .b(w234), .x(w861) );
	dmg_nand g786 (.a(w820), .b(w611), .x(w610) );
	dmg_nand g787 (.a(w188), .b(w824), .x(w821) );
	dmg_nand g788 (.a(w631), .b(w501), .x(w537) );
	dmg_nand g789 (.a(w400), .b(w401), .x(w411) );
	dmg_nand g790 (.a(w637), .b(w400), .x(w399) );
	dmg_nand g791 (.a(w1123), .b(w125), .x(w1148) );
	dmg_nand g792 (.a(w188), .b(w1297), .x(w915) );
	dmg_nand g793 (.a(w188), .b(w65), .x(w1178) );
	dmg_not2 g794 (.a(w1178), .x(w30) );
	dmg_nand g795 (.a(w637), .b(w1176), .x(w1177) );
	dmg_nand g796 (.a(w188), .b(w943), .x(w1006) );
	dmg_nand g797 (.a(w1131), .b(w611), .x(w67) );
	dmg_nand g798 (.a(w631), .b(w824), .x(w69) );
	dmg_nand g799 (.a(w997), .b(w933), .x(w1000) );
	dmg_nand g800 (.a(w637), .b(w829), .x(w828) );
	dmg_nand g801 (.a(w824), .b(w1091), .x(w1113) );
	dmg_nand g802 (.a(w824), .b(w1053), .x(w1052) );
	dmg_nand g803 (.a(w931), .b(w933), .x(w1077) );
	dmg_nand g804 (.a(w297), .b(w933), .x(w1187) );
	dmg_nand g805 (.a(w305), .b(w933), .x(w1306) );
	dmg_nand g806 (.a(w823), .b(w188), .x(w189) );
	dmg_nand g807 (.a(w331), .b(w294), .x(w304) );
	dmg_nand g808 (.a(w183), .b(w294), .x(w293) );
	dmg_nand g809 (.a(w943), .b(w1098), .x(w1101) );
	dmg_nand g810 (.a(w1035), .b(w188), .x(w1102) );
	dmg_nand g811 (.a(w631), .b(w943), .x(w944) );
	dmg_nand g812 (.a(w188), .b(w60), .x(w948) );
	dmg_nand g813 (.a(w412), .b(w60), .x(w413) );
	dmg_nand g814 (.a(w623), .b(w695), .x(w1206) );
	dmg_nand g815 (.a(w694), .b(w125), .x(w703) );
	dmg_nand g816 (.a(w693), .b(w125), .x(w1039) );
	dmg_nand g817 (.a(w188), .b(w637), .x(w709) );
	dmg_nand g818 (.a(w662), .b(w125), .x(w1249) );
	dmg_nand g819 (.a(w3), .b(w125), .x(w1145) );
	dmg_not6 g820 (.a(w387), .x(w388) );
	dmg_or g821 (.a(w90), .b(w1330), .x(w956) );
	dmg_or g822 (.a(w1087), .b(w231), .x(w1310) );
	dmg_or g823 (.a(w797), .b(w563), .x(w832) );
	dmg_or g824 (.a(w1068), .b(w1069), .x(w1065) );
	dmg_or g825 (.a(w70), .b(w340), .x(w979) );
	dmg_or g826 (.a(w614), .b(w615), .x(w1064) );
	dmg_or g827 (.a(w340), .b(w70), .x(w1181) );
	dmg_or g828 (.a(w1253), .b(w44), .x(w632) );
	dmg_or g829 (.a(w901), .b(w44), .x(w359) );
	dmg_or g830 (.a(w1208), .b(w93), .x(w94) );
	dmg_or g831 (.a(w1235), .b(w1130), .x(w774) );
	dmg_or g832 (.a(w772), .b(w469), .x(w424) );
	dmg_notif0 g833 (.n_ena(w225), .a(w1153), .x(w180) );
	dmg_notif0 g834 (.n_ena(w225), .a(w376), .x(w331) );
	dmg_notif0 g835 (.n_ena(w225), .a(w814), .x(w229) );
	dmg_notif0 g836 (.n_ena(w225), .a(w227), .x(w183) );
	dmg_notif0 g837 (.n_ena(w225), .a(w1151), .x(w16) );
	dmg_notif0 g838 (.n_ena(w225), .a(w1110), .x(w187) );
	dmg_notif0 g839 (.n_ena(w225), .a(w226), .x(w29) );
	dmg_notif0 g840 (.n_ena(w1052), .a(w987), .x(w183) );
	dmg_notif0 g841 (.n_ena(w310), .a(w940), .x(w183) );
	dmg_notif0 g842 (.n_ena(w310), .a(w1090), .x(w180) );
	dmg_notif0 g843 (.n_ena(w310), .a(w1080), .x(w331) );
	dmg_notif0 g844 (.n_ena(w310), .a(w941), .x(w55) );
	dmg_notif0 g845 (.n_ena(w310), .a(w1079), .x(w229) );
	dmg_notif0 g846 (.n_ena(w310), .a(w1076), .x(w29) );
	dmg_notif0 g847 (.n_ena(w310), .a(w309), .x(w16) );
	dmg_notif0 g848 (.n_ena(w15), .a(w20), .x(w183) );
	dmg_notif0 g849 (.n_ena(w15), .a(w20), .x(w16) );
	dmg_notif0 g850 (.n_ena(w15), .a(w20), .x(w180) );
	dmg_notif0 g851 (.n_ena(w15), .a(w20), .x(w229) );
	dmg_notif0 g852 (.n_ena(w15), .a(w20), .x(w331) );
	dmg_notif0 g853 (.n_ena(w15), .a(w20), .x(w55) );
	dmg_notif0 g854 (.n_ena(w643), .a(w35), .x(w55) );
	dmg_notif0 g855 (.n_ena(w643), .a(w36), .x(w187) );
	dmg_notif0 g856 (.n_ena(w413), .a(w630), .x(w187) );
	dmg_notif0 g857 (.n_ena(w993), .a(w994), .x(w180) );
	dmg_notif0 g858 (.n_ena(w993), .a(w1119), .x(w331) );
	dmg_notif0 g859 (.n_ena(w116), .a(w797), .x(w16) );
	dmg_notif0 g860 (.n_ena(w812), .a(w1093), .x(w29) );
	dmg_notif0 g861 (.n_ena(w812), .a(w840), .x(w55) );
	dmg_notif0 g862 (.n_ena(w828), .a(w827), .x(w183) );
	dmg_notif0 g863 (.n_ena(w812), .a(w1049), .x(w187) );
	dmg_notif0 g864 (.n_ena(w812), .a(w1073), .x(w16) );
	dmg_notif0 g865 (.n_ena(w1113), .a(w77), .x(w55) );
	dmg_notif0 g866 (.n_ena(w812), .a(w817), .x(w180) );
	dmg_notif0 g867 (.n_ena(w812), .a(w1105), .x(w331) );
	dmg_notif0 g868 (.n_ena(w1177), .a(w965), .x(w331) );
	dmg_notif0 g869 (.n_ena(w548), .a(w739), .x(w55) );
	dmg_notif0 g870 (.n_ena(w526), .a(w1321), .x(w16) );
	dmg_notif0 g871 (.n_ena(w526), .a(w1323), .x(w29) );
	dmg_notif0 g872 (.n_ena(w526), .a(w525), .x(w187) );
	dmg_notif0 g873 (.n_ena(w359), .a(w358), .x(w229) );
	dmg_notif0 g874 (.n_ena(w411), .a(w410), .x(w187) );
	dmg_notif0 g875 (.n_ena(w505), .a(w506), .x(w55) );
	dmg_notif0 g876 (.n_ena(w28), .a(w1191), .x(w55) );
	dmg_notif0 g877 (.n_ena(w28), .a(w535), .x(w16) );
	dmg_notif0 g878 (.n_ena(w28), .a(w329), .x(w331) );
	dmg_notif0 g879 (.n_ena(w474), .a(w971), .x(w29) );
	dmg_notif0 g880 (.n_ena(w474), .a(w1111), .x(w55) );
	dmg_notif0 g881 (.n_ena(w474), .a(w972), .x(w16) );
	dmg_notif0 g882 (.n_ena(w483), .a(w1370), .x(w16) );
	dmg_notif0 g883 (.n_ena(w483), .a(w616), .x(w229) );
	dmg_notif0 g884 (.n_ena(w116), .a(w779), .x(w229) );
	dmg_notif0 g885 (.n_ena(w432), .a(w431), .x(w187) );
	dmg_notif0 g886 (.n_ena(w212), .a(w1283), .x(w331) );
	dmg_notif0 g887 (.n_ena(w212), .a(w1228), .x(w183) );
	dmg_notif0 g888 (.n_ena(w212), .a(w374), .x(w180) );
	dmg_notif0 g889 (.n_ena(w177), .a(w462), .x(w229) );
	dmg_notif0 g890 (.n_ena(w177), .a(w634), .x(w183) );
	dmg_notif0 g891 (.n_ena(w177), .a(w636), .x(w16) );
	dmg_notif0 g892 (.n_ena(w609), .a(w1351), .x(w331) );
	dmg_notif0 g893 (.n_ena(w609), .a(w608), .x(w180) );
	dmg_notif0 g894 (.n_ena(w177), .a(w192), .x(w29) );
	dmg_notif0 g895 (.n_ena(w174), .a(w1287), .x(w331) );
	dmg_notif0 g896 (.n_ena(w174), .a(w184), .x(w183) );
	dmg_notif0 g897 (.n_ena(w177), .a(w186), .x(w187) );
	dmg_notif0 g898 (.n_ena(w177), .a(w459), .x(w55) );
	dmg_notif0 g899 (.n_ena(w177), .a(w447), .x(w331) );
	dmg_notif0 g900 (.n_ena(w177), .a(w178), .x(w180) );
	dmg_notif0 g901 (.n_ena(w116), .a(w620), .x(w29) );
	dmg_notif0 g902 (.n_ena(w28), .a(w1128), .x(w29) );
	dmg_notif0 g903 (.n_ena(w28), .a(w256), .x(w229) );
	dmg_notif0 g904 (.n_ena(w28), .a(w569), .x(w180) );
	dmg_notif0 g905 (.n_ena(w116), .a(w776), .x(w183) );
	dmg_notif0 g906 (.n_ena(w116), .a(w117), .x(w180) );
	dmg_notif0 g907 (.n_ena(w909), .a(w782), .x(w229) );
	dmg_notif0 g908 (.n_ena(w46), .a(w138), .x(w183) );
	dmg_notif0 g909 (.n_ena(w46), .a(w332), .x(w331) );
	dmg_notif0 g910 (.n_ena(w46), .a(w1272), .x(w180) );
	dmg_notif0 g911 (.n_ena(w47), .a(w1012), .x(w229) );
	dmg_notif0 g912 (.n_ena(w483), .a(w54), .x(w55) );
	dmg_notif0 g913 (.n_ena(w483), .a(w482), .x(w187) );
	dmg_notif0 g914 (.n_ena(w483), .a(w1270), .x(w29) );
	dmg_notif0 g915 (.n_ena(w474), .a(w475), .x(w187) );
	dmg_notif0 g916 (.n_ena(w432), .a(w433), .x(w229) );
	dmg_notif0 g917 (.n_ena(w432), .a(w849), .x(w55) );
	dmg_notif0 g918 (.n_ena(w432), .a(w850), .x(w29) );
	dmg_notif0 g919 (.n_ena(w499), .a(w498), .x(w55) );
	dmg_notif0 g920 (.n_ena(w432), .a(w213), .x(w16) );
	dmg_notif0 g921 (.n_ena(w1254), .a(w1235), .x(w187) );
	dmg_notif0 g922 (.n_ena(w359), .a(w350), .x(w16) );
	dmg_notif0 g923 (.n_ena(w359), .a(w349), .x(w55) );
	dmg_notif0 g924 (.n_ena(w359), .a(w557), .x(w29) );
	dmg_notif0 g925 (.n_ena(w359), .a(w360), .x(w187) );
	dmg_notif0 g926 (.n_ena(w632), .a(w729), .x(w183) );
	dmg_notif0 g927 (.n_ena(w632), .a(w364), .x(w331) );
	dmg_notif0 g928 (.n_ena(w632), .a(w633), .x(w180) );
	dmg_notif0 g929 (.n_ena(w907), .a(w588), .x(w16) );
	dmg_notif0 g930 (.n_ena(w907), .a(w590), .x(w55) );
	dmg_notif0 g931 (.n_ena(w609), .a(w908), .x(w183) );
	dmg_notif0 g932 (.n_ena(w174), .a(w1258), .x(w180) );
	dmg_notif0 g933 (.n_ena(w555), .a(w1262), .x(w183) );
	dmg_notif0 g934 (.n_ena(w555), .a(w654), .x(w29) );
	dmg_notif0 g935 (.n_ena(w555), .a(w669), .x(w331) );
	dmg_notif0 g936 (.n_ena(w555), .a(w107), .x(w180) );
	dmg_notif0 g937 (.n_ena(w548), .a(w747), .x(w183) );
	dmg_notif0 g938 (.n_ena(w555), .a(w106), .x(w229) );
	dmg_notif0 g939 (.n_ena(w548), .a(w1212), .x(w229) );
	dmg_notif0 g940 (.n_ena(w548), .a(w740), .x(w331) );
	dmg_notif0 g941 (.n_ena(w548), .a(w1240), .x(w180) );
	dmg_notif0 g942 (.n_ena(w399), .a(w398), .x(w180) );
	dmg_notif0 g943 (.n_ena(w28), .a(w912), .x(w187) );
	dmg_notif0 g944 (.n_ena(w28), .a(w326), .x(w183) );
	dmg_notif0 g945 (.n_ena(w68), .a(w1005), .x(w331) );
	dmg_notif0 g946 (.n_ena(w68), .a(w825), .x(w180) );
	dmg_notif0 g947 (.n_ena(w68), .a(w911), .x(w183) );
	dmg_notif0 g948 (.n_ena(w993), .a(w967), .x(w183) );
	dmg_notif0 g949 (.n_ena(w413), .a(w484), .x(w55) );
	dmg_notif0 g950 (.n_ena(w1101), .a(w1100), .x(w55) );
	dmg_notif0 g951 (.n_ena(w15), .a(w20), .x(w29) );
	dmg_notif0 g952 (.n_ena(w15), .a(w20), .x(w187) );
	dmg_notif0 g953 (.n_ena(w812), .a(w1154), .x(w183) );
	dmg_notif0 g954 (.n_ena(w812), .a(w813), .x(w229) );
	dmg_notif0 g955 (.n_ena(w225), .a(w224), .x(w55) );
	dmg_and g956 (.a(w1061), .b(w132), .x(w131) );
	dmg_and g957 (.a(w133), .b(w132), .x(w1071) );
	dmg_and g958 (.a(w933), .b(w1313), .x(w1312) );
	dmg_and g959 (.a(w933), .b(w1044), .x(w1045) );
	dmg_and g960 (.a(w156), .b(w155), .x(w545) );
	dmg_and g961 (.a(w440), .b(w155), .x(w544) );
	dmg_and g962 (.a(w541), .b(w155), .x(w543) );
	dmg_and g963 (.a(w471), .b(w155), .x(w542) );
	dmg_and g964 (.a(w294), .b(w547), .x(w546) );
	dmg_and g965 (.a(w294), .b(w1347), .x(w1346) );
	dmg_and g966 (.a(w355), .b(w354), .x(w1345) );
	dmg_and g967 (.a(w1209), .b(w354), .x(w1344) );
	dmg_and g968 (.a(w353), .b(w354), .x(w1343) );
	dmg_and g969 (.a(w91), .b(w354), .x(w1328) );
	dmg_and g970 (.a(w1202), .b(w188), .x(w631) );
	dmg_and g971 (.a(w1342), .b(w880), .x(w801) );
	dmg_and g972 (.a(w713), .b(w798), .x(w1038) );
	dmg_and g973 (.a(w188), .b(w60), .x(w624) );
	dmg_and g974 (.a(w924), .b(w925), .x(w1266) );
	dmg_and g975 (.a(w24), .b(w23), .x(w22) );
	dmg_and g976 (.a(w826), .b(w914), .x(w154) );
	dmg_and g977 (.a(w188), .b(w313), .x(w142) );
	dmg_and g978 (.a(w831), .b(w830), .x(w1053) );
	dmg_and g979 (.a(w838), .b(w271), .x(w986) );
	dmg_and g980 (.a(w223), .b(w611), .x(w612) );
	dmg_and g981 (.a(w76), .b(w75), .x(w1070) );
	dmg_and g982 (.a(w236), .b(w873), .x(w869) );
	dmg_and g983 (.a(w236), .b(w966), .x(w1116) );
	dmg_and g984 (.a(w30), .b(w763), .x(w762) );
	dmg_and g985 (.a(w30), .b(w512), .x(w761) );
	dmg_and g986 (.a(w487), .b(w488), .x(w493) );
	dmg_and g987 (.a(w493), .b(w492), .x(w627) );
	dmg_and g988 (.a(w30), .b(w31), .x(w1324) );
	dmg_and g989 (.a(w317), .b(w316), .x(w42) );
	dmg_and g990 (.a(w32), .b(w895), .x(w896) );
	dmg_and g991 (.a(w902), .b(w188), .x(w1211) );
	dmg_and g992 (.a(w904), .b(w188), .x(w1251) );
	dmg_and g993 (.a(w29), .b(w90), .x(w1252) );
	dmg_and g994 (.a(w188), .b(w637), .x(w638) );
	dmg_and g995 (.a(w188), .b(w902), .x(w674) );
	dmg_and g996 (.a(w496), .b(w497), .x(w1195) );
	dmg_and g997 (.a(w401), .b(w188), .x(w1194) );
	dmg_and g998 (.a(w210), .b(w188), .x(w1282) );
	dmg_and g999 (.a(w886), .b(w188), .x(w810) );
	dmg_and g1000 (.a(w188), .b(w42), .x(w975) );
	dmg_and g1001 (.a(w1011), .b(w478), .x(w1010) );
	dmg_and g1002 (.a(w234), .b(w790), .x(w791) );
	dmg_and g1003 (.a(w234), .b(w792), .x(w1379) );
	dmg_and g1004 (.a(w452), .b(w188), .x(w200) );
	dmg_and g1005 (.a(w504), .b(w188), .x(w451) );
	dmg_and g1006 (.a(w452), .b(w188), .x(w203) );
	dmg_and g1007 (.a(w30), .b(w466), .x(w1274) );
	dmg_and g1008 (.a(w30), .b(w1232), .x(w1127) );
	dmg_and g1009 (.a(w234), .b(w270), .x(w250) );
	dmg_and g1010 (.a(w236), .b(w865), .x(w238) );
	dmg_and g1011 (.a(w236), .b(w237), .x(w240) );
	dmg_and g1012 (.a(w188), .b(w42), .x(w1271) );
	dmg_and g1013 (.a(w188), .b(w210), .x(w724) );
	dmg_and g1014 (.a(w188), .b(w454), .x(w1355) );
	dmg_and g1015 (.a(w501), .b(w188), .x(w181) );
	dmg_and g1016 (.a(w1259), .b(w686), .x(w597) );
	dmg_and g1017 (.a(w658), .b(w659), .x(w655) );
	dmg_and g1018 (.a(w1241), .b(w1242), .x(w670) );
	dmg_and g1019 (.a(w30), .b(w527), .x(w528) );
	dmg_and g1020 (.a(w30), .b(w1184), .x(w976) );
	dmg_and g1021 (.a(w30), .b(w327), .x(w328) );
	dmg_and g1022 (.a(w76), .b(w611), .x(w831) );
	dmg_and g1023 (.a(w166), .b(w162), .x(w163) );
	dmg_and g1024 (.a(w188), .b(w943), .x(w294) );
	dmg_and g1025 (.a(w188), .b(w886), .x(w1179) );
	dmg_and g1026 (.a(w760), .b(w508), .x(w507) );
	dmg_and g1027 (.a(w889), .b(w892), .x(w32) );
	dmg_and g1028 (.a(w317), .b(w318), .x(w637) );
	dmg_and g1029 (.a(w586), .b(w524), .x(w715) );
	dmg_and g1030 (.a(w397), .b(w647), .x(w754) );
	dmg_and g1031 (.a(w397), .b(w716), .x(w1334) );
	dmg_and g1032 (.a(w397), .b(w717), .x(w1037) );
	dmg_and g1033 (.a(w397), .b(w715), .x(w714) );
	dmg_and g1034 (.a(w188), .b(w204), .x(w1122) );
	dmg_and g1035 (.a(w188), .b(w695), .x(w574) );
	dmg_and g1036 (.a(w294), .b(w1348), .x(w1349) );
	dmg_and g1037 (.a(w933), .b(w998), .x(w1314) );
	dmg_and g1038 (.a(w1088), .b(w1089), .x(w258) );
	dmg_and g1039 (.a(w129), .b(w132), .x(w130) );
	dmg_and g1040 (.a(w834), .b(w132), .x(w1152) );
	dmg_nand4 g1041 (.a(w1204), .b(w1200), .c(w578), .d(w111), .x(w1201) );
	dmg_nand4 g1042 (.a(w951), .b(w113), .c(w800), .d(w801), .x(w570) );
	dmg_nand4 g1043 (.a(w207), .b(w62), .c(w315), .d(w640), .x(w639) );
	dmg_nand4 g1044 (.a(w208), .b(w315), .c(w62), .d(w209), .x(w991) );
	dmg_nand4 g1045 (.a(w209), .b(w63), .c(w315), .d(w640), .x(w503) );
	dmg_nand4 g1046 (.a(w640), .b(w206), .c(w63), .d(w209), .x(w641) );
	dmg_nand4 g1047 (.a(w207), .b(w63), .c(w206), .d(w640), .x(w642) );
	dmg_nand4 g1048 (.a(w208), .b(w206), .c(w63), .d(w207), .x(w64) );
	dmg_nand4 g1049 (.a(w209), .b(w62), .c(w315), .d(w640), .x(w720) );
	dmg_nand4 g1050 (.a(w209), .b(w62), .c(w315), .d(w208), .x(w1036) );
	dmg_nand4 g1051 (.a(w208), .b(w206), .c(w62), .d(w209), .x(w314) );
	dmg_nand4 g1052 (.a(w208), .b(w206), .c(w63), .d(w209), .x(w402) );
	dmg_nand4 g1053 (.a(w208), .b(w315), .c(w63), .d(w209), .x(w205) );
	dmg_nand4 g1054 (.a(w207), .b(w63), .c(w206), .d(w208), .x(w1041) );
	dmg_nand4 g1055 (.a(w640), .b(w206), .c(w62), .d(w207), .x(w1149) );
	dmg_nand4 g1056 (.a(w207), .b(w62), .c(w206), .d(w208), .x(w1248) );
	dmg_nand4 g1057 (.a(w208), .b(w206), .c(w62), .d(w207), .x(w61) );
	dmg_nand4 g1058 (.a(w207), .b(w62), .c(w315), .d(w208), .x(w990) );
	dmg_nand4 g1059 (.a(w208), .b(w315), .c(w63), .d(w207), .x(w903) );
	dmg_nand4 g1060 (.a(w640), .b(w206), .c(w62), .d(w209), .x(w1173) );
	dmg_nand4 g1061 (.a(w209), .b(w62), .c(w206), .d(w208), .x(w962) );
	dmg_mux g1062 (.sel(w397), .d1(w102), .d0(w103), .q(w1340) );
	dmg_mux g1063 (.sel(w397), .d1(w105), .d0(w104), .q(w1142) );
	dmg_mux g1064 (.sel(w397), .d1(w109), .d0(w110), .q(w1143) );
	dmg_mux g1065 (.sel(w397), .d1(w396), .d0(w707), .q(w1164) );
	dmg_mux g1066 (.sel(w383), .d1(w381), .d0(w382), .q(w1331) );
	dmg_mux g1067 (.sel(w383), .d1(w576), .d0(w577), .q(w1237) );
	dmg_mux g1068 (.sel(w383), .d1(w1341), .d0(w4), .q(w3) );
	dmg_mux g1069 (.sel(w383), .d1(w1125), .d0(w1124), .q(w662) );
	dmg_mux g1070 (.sel(w383), .d1(w385), .d0(w384), .q(w1123) );
	dmg_mux g1071 (.sel(w383), .d1(w691), .d0(w692), .q(w693) );
	dmg_mux g1072 (.sel(w383), .d1(w579), .d0(w690), .q(w694) );
	dmg_mux g1073 (.sel(w383), .d1(w7), .d0(w6), .q(w128) );
	dmg_mux g1074 (.sel(w831), .d1(w476), .d0(w1010), .q(w613) );
	dmg_mux g1075 (.sel(w1029), .d1(w141), .d0(w263), .q(w858) );
	dmg_mux g1076 (.sel(w973), .d1(w1066), .d0(w1065), .q(w476) );
	dmg_mux g1077 (.sel(w1029), .d1(w141), .d0(w1188), .q(w1305) );
	dmg_mux g1078 (.sel(w1029), .d1(w141), .d0(w1042), .q(w1296) );
	dmg_mux g1079 (.sel(w397), .d1(w379), .d0(w582), .q(w1332) );
	dmg_mux g1080 (.sel(w397), .d1(w668), .d0(w667), .q(w1141) );
	dmg_bufif0 g1081 (.a0(w1146), .n_ena(w125), .a1(w1146), .x(w104) );
	dmg_bufif0 g1082 (.a0(w124), .n_ena(w125), .a1(w124), .x(w111) );
	dmg_bufif0 g1083 (.a0(w689), .n_ena(w125), .a1(w689), .x(w110) );
	dmg_bufif0 g1084 (.a0(w1161), .n_ena(w125), .a1(w1161), .x(w578) );
	dmg_bufif0 g1085 (.a0(w87), .n_ena(w125), .a1(w87), .x(w666) );
	dmg_bufif0 g1086 (.a0(w989), .n_ena(w125), .a1(w989), .x(w112) );
	dmg_bufif0 g1087 (.a0(w699), .n_ena(w125), .a1(w699), .x(w103) );
	dmg_nor_latch g1088 (.s(w733), .r(w683), .q(w682) );
	dmg_nor_latch g1089 (.s(w565), .r(w426), .q(w427) );
	dmg_nor_latch g1090 (.s(w854), .r(w120), .nq(w855) );
	dmg_nor_latch g1091 (.s(w340), .r(w837), .q(w1011) );
	dmg_nor_latch g1092 (.s(w1267), .r(w979), .q(w978) );
	dmg_nor_latch g1093 (.s(w917), .r(w920), .nq(w919) );
	dmg_nor_latch g1094 (.s(w346), .r(w407), .q(w406) );
	dmg_nor_latch g1095 (.s(w738), .r(w595), .nq(w737) );
	dmg_nor_latch g1096 (.s(w745), .r(w742), .nq(w743) );
	dmg_nor_latch g1097 (.s(w347), .r(w923), .q(w924) );
	dmg_nor_latch g1098 (.s(w27), .r(w1303), .q(w826) );
	dmg_bufif0 g1099 (.a0(w443), .n_ena(w125), .a1(w443), .x(w667) );
	dmg_not2 g1100 (.a(w395), .x(w396) );
	dmg_latch g1101 (.ena(w5), .d(w103), .q(w382) );
	dmg_latch g1102 (.ena(w5), .d(w578), .q(w4) );
	dmg_latch g1103 (.ena(w5), .d(w112), .q(w577) );
	dmg_latch g1104 (.ena(w5), .d(w110), .q(w1124) );
	dmg_latch g1105 (.ena(w5), .d(w666), .q(w384) );
	dmg_latch g1106 (.ena(w5), .d(w111), .q(w690) );
	dmg_latch g1107 (.ena(w5), .d(w667), .q(w6) );
	dmg_latch g1108 (.ena(w5), .d(w104), .q(w692) );
	dmg_latch g1109 (.ena(w10), .d(w879), .q(w1203) );
	dmg_latch g1110 (.ena(w116), .d(w781), .q(w117) );
	dmg_latch g1111 (.ena(w116), .d(w777), .q(w776) );
	dmg_latch g1112 (.ena(w116), .d(w778), .q(w436) );
	dmg_latch g1113 (.ena(w116), .d(w780), .q(w779) );
	dmg_not4 g1114 (.a(w143), .x(w144) );
	dmg_dffsr g1115 (.nset1(w1077), .nset2(w1077), .d(w306), .q(w1078), .nres(w1311), .clk(w1043) );
	dmg_dffsr g1116 (.nset1(w304), .nset2(w304), .d(w1032), .q(w931), .nres(w1183), .clk(w1033) );
	dmg_dffsr g1117 (.nset1(w884), .nset2(w884), .d(w883), .q(w566), .nres(w1374), .clk(w258) );
	dmg_dffsr g1118 (.nset1(w1000), .nset2(w1000), .d(w1001), .q(w301), .nres(w999), .clk(w1043) );
	dmg_dffsr g1119 (.nset1(w1187), .nset2(w1187), .d(w1078), .q(w1001), .nres(w1327), .clk(w1043) );
	dmg_dffsr g1120 (.nset1(w1371), .nset2(w1371), .d(w794), .q(w793), .nres(w864), .clk(w219) );
	dmg_dffsr g1121 (.nset1(w259), .nset2(w259), .d(w805), .q(w789), .nres(w215), .clk(w258) );
	dmg_dffsr g1122 (.nset1(w253), .nset2(w253), .d(w871), .q(w232), .nres(w216), .clk(w217) );
	dmg_dffsr g1123 (.nset1(w796), .nset2(w796), .d(w232), .q(w794), .nres(w239), .clk(w217) );
	dmg_dffsr g1124 (.nset1(w235), .nset2(w235), .d(w793), .q(w862), .nres(w785), .clk(w219) );
	dmg_dffsr g1125 (.nset1(w558), .nset2(w558), .d(w1216), .q(w764), .nres(w1214), .clk(w258) );
	dmg_dffsr g1126 (.nset1(w172), .nset2(w172), .d(w1129), .q(w997), .nres(w1325), .clk(w258) );
	dmg_dffsr g1127 (.nset1(w788), .nset2(w788), .d(w787), .q(w567), .nres(w472), .clk(w258) );
	dmg_dffsr g1128 (.nset1(w1326), .nset2(w1326), .d(w769), .q(w874), .nres(w936), .clk(w258) );
	dmg_dffsr g1129 (.nset1(w1114), .nset2(w1114), .d(w415), .q(w860), .nres(w414), .clk(w258) );
	dmg_dffsr g1130 (.nset1(w861), .nset2(w861), .d(w862), .q(w268), .nres(w269), .clk(w219) );
	dmg_dffsr g1131 (.nset1(w264), .nset2(w264), .d(w265), .q(w871), .nres(w870), .clk(w217) );
	dmg_dffsr g1132 (.nset1(w302), .nset2(w302), .d(w301), .q(w265), .nres(w1185), .clk(w217) );
	dmg_dffsr g1133 (.nset1(w417), .nset2(w417), .d(w419), .q(w254), .nres(w418), .clk(w258) );
	dmg_dffsr g1134 (.nset1(w293), .nset2(w293), .d(w1004), .q(w297), .nres(w296), .clk(w1033) );
	dmg_dffsr g1135 (.nset1(w1306), .nset2(w1306), .d(w20), .q(w306), .nres(w1315), .clk(w1043) );
	dmg_not6 g1136 (.a(w44), .x(w623) );
	dmg_not6 g1137 (.a(w706), .x(w707) );
	dmg_mux g1138 (.sel(w611), .d1(w85), .d0(w957), .q(w84) );
	dmg_not6 g1139 (.a(w799), .x(w188) );
	dmg_not6 g1140 (.a(w1210), .x(w611) );
	dmg_not6 g1141 (.a(w775), .x(w70) );
	dmg_dffr_comp g1142 (.nr1(w298), .nr2(w298), .d(w266), .ck(w144), .cck(w773), .q(w252) );
	dmg_dffr_comp g1143 (.nr1(w298), .nr2(w298), .d(w789), .ck(w144), .cck(w468), .q(w423) );
	dmg_dffr_comp g1144 (.nr1(w298), .nr2(w298), .d(w875), .ck(w144), .cck(w768), .q(w1389) );
	dmg_dffr_comp g1145 (.nr1(w298), .nr2(w298), .d(w566), .ck(w144), .cck(w468), .q(w251) );
	dmg_dffr_comp g1146 (.nr1(w298), .nr2(w298), .d(w254), .ck(w144), .cck(w765), .q(w771) );
	dmg_dffr_comp g1147 (.nr1(w298), .nr2(w298), .d(w860), .ck(w144), .cck(w468), .q(w934) );
	dmg_dffr_comp g1148 (.nr1(w298), .nr2(w298), .d(w416), .ck(w144), .cck(w768), .q(w767) );
	dmg_dffr_comp g1149 (.nr1(w298), .nr2(w298), .d(w868), .ck(w144), .cck(w299), .q(w866) );
	dmg_dffr_comp g1150 (.nr1(w298), .nr2(w298), .d(w935), .ck(w144), .cck(w299), .q(w872) );
	dmg_dffr_comp g1151 (.nr1(w298), .nr2(w298), .d(w300), .ck(w144), .cck(w299), .q(w928) );
	dmg_dffr_comp g1152 (.nr1(w298), .nr2(w298), .d(w764), .ck(w144), .cck(w930), .q(w1030) );
	dmg_dffr_comp g1153 (.nr1(w298), .nr2(w298), .d(w1132), .ck(w144), .cck(w299), .q(w927) );
	dmg_dffr_comp g1154 (.nr1(w298), .nr2(w298), .d(w931), .ck(w144), .cck(w930), .q(w867) );
	dmg_dffr_comp g1155 (.nr1(w298), .nr2(w298), .d(w267), .ck(w144), .cck(w773), .q(w807) );
	dmg_dffr_comp g1156 (.nr1(w298), .nr2(w298), .d(w863), .ck(w144), .cck(w773), .q(w786) );
	dmg_dffr_comp g1157 (.nr1(w298), .nr2(w298), .d(w859), .ck(w144), .cck(w773), .q(w795) );
	dmg_dffr_comp g1158 (.nr1(w298), .nr2(w298), .d(w567), .ck(w144), .cck(w468), .q(w467) );
	dmg_dffr_comp g1159 (.nr1(w298), .nr2(w298), .d(w305), .ck(w144), .cck(w765), .q(w1386) );
	dmg_dffr_comp g1160 (.nr1(w298), .nr2(w298), .d(w997), .ck(w144), .cck(w930), .q(w929) );
	dmg_dffr_comp g1161 (.nr1(w298), .nr2(w298), .d(w1002), .ck(w144), .cck(w768), .q(w1385) );
	dmg_dffr_comp g1162 (.nr1(w298), .nr2(w298), .d(w297), .ck(w144), .cck(w930), .q(w926) );
	dmg_not4 g1163 (.a(w123), .x(w122) );
	dmg_dffr_comp g1164 (.nr1(w298), .nr2(w298), .d(w874), .ck(w144), .cck(w765), .q(w766) );
	dmg_or g1165 (.a(w45), .b(w44), .x(w46) );
	dmg_or g1166 (.a(w43), .b(w44), .x(w474) );
	dmg_or g1167 (.a(w1362), .b(w1363), .x(w48) );
	dmg_or g1168 (.a(w70), .b(w27), .x(w437) );
	dmg_or g1169 (.a(w70), .b(w27), .x(w426) );
	dmg_or g1170 (.a(w620), .b(w563), .x(w562) );
	dmg_or g1171 (.a(w1220), .b(w44), .x(w432) );
	dmg_or g1172 (.a(w211), .b(w44), .x(w212) );
	dmg_or g1173 (.a(w721), .b(w610), .x(w609) );
	dmg_or g1174 (.a(w70), .b(w347), .x(w683) );
	dmg_or g1175 (.a(w1339), .b(w175), .x(w174) );
	dmg_or g1176 (.a(w992), .b(w67), .x(w68) );
	dmg_or g1177 (.a(w613), .b(w612), .x(w132) );
	dmg_or g1178 (.a(w154), .b(w611), .x(w155) );
	dmg_or g1179 (.a(w1266), .b(w611), .x(w354) );
	dmg_or g1180 (.a(w1099), .b(w44), .x(w993) );
	dmg_or g1181 (.a(w1197), .b(w1198), .x(w887) );
	dmg_aon22 g1182 (.a0(w134), .a1(w1061), .b0(w1268), .b1(w616), .x(w1062) );
	dmg_aon22 g1183 (.a0(w134), .a1(w129), .b0(w1060), .b1(w616), .x(w1063) );
	dmg_aon22 g1184 (.a0(w134), .a1(w133), .b0(w980), .b1(w616), .x(w835) );
	dmg_aon22 g1185 (.a0(w502), .a1(w673), .b0(w673), .b1(w358), .x(w900) );
	dmg_aon22 g1186 (.a0(w502), .a1(w353), .b0(w899), .b1(w358), .x(w898) );
	dmg_aon22 g1187 (.a0(w502), .a1(w91), .b0(w897), .b1(w358), .x(w357) );
	dmg_aon22 g1188 (.a0(w502), .a1(w355), .b0(w356), .b1(w358), .x(w362) );
	dmg_aon22 g1189 (.a0(w648), .a1(w524), .b0(w586), .b1(w649), .x(w717) );
	dmg_aon22 g1190 (.a0(w439), .a1(w440), .b0(w441), .b1(w433), .x(w531) );
	dmg_aon22 g1191 (.a0(w439), .a1(w434), .b0(w434), .b1(w433), .x(w442) );
	dmg_aon22 g1192 (.a0(w439), .a1(w541), .b0(w533), .b1(w433), .x(w847) );
	dmg_aon22 g1193 (.a0(w439), .a1(w156), .b0(w532), .b1(w433), .x(w157) );
	dmg_aon22 g1194 (.a0(w51), .a1(w783), .b0(w782), .b1(w784), .x(w246) );
	dmg_muxi g1195 (.sel(w521), .d1(w518), .d0(w517), .q(w648) );
	dmg_muxi g1196 (.sel(w521), .d1(w520), .d0(w585), .q(w586) );
	dmg_muxi g1197 (.sel(w618), .d1(w56), .d0(w57), .q(w1233) );
	dmg_muxi g1198 (.sel(w521), .d1(w522), .d0(w1247), .q(w523) );
	dmg_muxi g1199 (.sel(w521), .d1(w751), .d0(w752), .q(w718) );
	dmg_nand_latch g1200 (.nr(w344), .ns(w684), .nq(w685) );
	dmg_nand_latch g1201 (.nr(w145), .ns(w150), .nq(w146) );
	dmg_nand_latch g1202 (.nr(w1361), .ns(w1360), .nq(w1362) );
	dmg_nand_latch g1203 (.nr(w959), .ns(w98), .nq(w99) );
	dmg_not g1204 (.a(w553), .x(w554) );
	dmg_nand g1205 (.a(w1121), .b(w204), .x(w643) );
	dmg_nand g1206 (.a(w188), .b(w504), .x(w1172) );
	dmg_nand g1207 (.a(w42), .b(w188), .x(w334) );
	dmg_nor3 g1208 (.a(w1016), .b(w983), .c(w982), .x(w1017) );
	dmg_nor3 g1209 (.a(w1016), .b(w972), .c(w982), .x(w984) );
	dmg_nor3 g1210 (.a(w1016), .b(w983), .c(w971), .x(w1019) );
	dmg_nor3 g1211 (.a(w1111), .b(w983), .c(w982), .x(w221) );
	dmg_nor3 g1212 (.a(w1111), .b(w972), .c(w971), .x(w273) );
	dmg_nor3 g1213 (.a(w1111), .b(w972), .c(w982), .x(w981) );
	dmg_nor3 g1214 (.a(w75), .b(w1008), .c(w77), .x(w78) );
	dmg_nor3 g1215 (.a(w1111), .b(w983), .c(w971), .x(w842) );
	dmg_nor3 g1216 (.a(w70), .b(w27), .c(w163), .x(w164) );
	dmg_nor3 g1217 (.a(w760), .b(w1008), .c(w506), .x(w1175) );
	dmg_nor3 g1218 (.a(w947), .b(w70), .c(w27), .x(w26) );
	dmg_nor3 g1219 (.a(w24), .b(w1008), .c(w1100), .x(w1293) );
	dmg_nor3 g1220 (.a(w1016), .b(w972), .c(w971), .x(w970) );
	dmg_nor3 g1221 (.a(w72), .b(w70), .c(w340), .x(w73) );
	dmg_nor3 g1222 (.a(w1117), .b(w1118), .c(w1182), .x(w977) );
	dmg_nor3 g1223 (.a(w496), .b(w1008), .c(w498), .x(w1281) );
	dmg_nor3 g1224 (.a(w1285), .b(w1284), .c(w429), .x(w428) );
	dmg_nor3 g1225 (.a(w1219), .b(w70), .c(w346), .x(w539) );
	dmg_nor3 g1226 (.a(w728), .b(w1257), .c(w1256), .x(w681) );
	dmg_nor3 g1227 (.a(w70), .b(w347), .c(w670), .x(w671) );
	dmg_nor3 g1228 (.a(w70), .b(w346), .c(w597), .x(w596) );
	dmg_nor3 g1229 (.a(w70), .b(w346), .c(w655), .x(w656) );
	dmg_nand_latch g1230 (.nr(w322), .ns(w885), .nq(w323) );
	dmg_nand g1231 (.a(w188), .b(w1218), .x(w320) );
	dmg_not g1232 (.a(w305), .x(w1313) );
	dmg_dffsr g1233 (.nset1(w1309), .nset2(w1309), .d(w1085), .q(w305), .nres(w1308), .clk(w1033) );
	dmg_not6 g1234 (.a(w114), .x(w44) );
	dmg_nor3 g1235 (.a(w1159), .b(w70), .c(w347), .x(w1169) );
	dmg_fa g1236 (.cin(w422), .s(w787), .cout(w421), .a(w467), .b(w786) );
	dmg_fa g1237 (.cin(w421), .s(w883), .cout(w420), .a(w251), .b(w252) );
	dmg_fa g1238 (.cin(w231), .s(w415), .cout(w806), .a(w934), .b(w807) );
	dmg_fa g1239 (.cin(w770), .s(w769), .cout(w1387), .a(w766), .b(w767) );
	dmg_fa g1240 (.cin(w1215), .s(w1129), .cout(w1003), .a(w929), .b(w928) );
	dmg_fa g1241 (.cin(w1387), .s(w1216), .cout(w1215), .a(w1030), .b(w872) );
	dmg_fa g1242 (.cin(w806), .s(w805), .cout(w422), .a(w423), .b(w795) );
	dmg_fa g1243 (.cin(w420), .s(w419), .cout(w770), .a(w771), .b(w1389) );
	dmg_fa g1244 (.cin(w1186), .s(w1032), .cout(w1031), .a(w867), .b(w866) );
	dmg_fa g1245 (.cin(w1003), .s(w1004), .cout(w1186), .a(w926), .b(w927) );
	dmg_fa g1246 (.cin(w1031), .s(w1085), .cout(w1086), .a(w1386), .b(w1385) );
	dmg_aon222 g1247 (.a0(w523), .a1(w524), .b0(w718), .b1(w649), .c0(w648), .c1(w587), .x(w647) );
	dmg_aon222 g1248 (.a0(w718), .a1(w524), .b0(w648), .b1(w649), .c0(w586), .c1(w587), .x(w716) );
	dmg_aon22 g1249 (.a0(w134), .a1(w135), .b0(w135), .b1(w616), .x(w617) );
	dmg_aon222222 g1250 (.a0(w843), .a1(w842), .b0(w220), .b1(w221), .c0(w277), .c1(w970), .d0(w1009), .d1(w984), .e0(w276), .e1(w1019), .f0(w1021), .f1(w1017), .x(w1066) );
	dmg_aon2222 g1251 (.a0(w274), .a1(w273), .b0(w272), .b1(w981), .c0(w841), .c1(w842), .d0(w222), .d1(w221), .x(w1069) );
	dmg_aon2222 g1252 (.a0(w1054), .a1(w970), .b0(w985), .b1(w984), .c0(w1015), .c1(w1019), .d0(w1018), .d1(w1017), .x(w1068) );
	dmg_aon2222 g1253 (.a0(w627), .a1(w628), .b0(w493), .b1(w1301), .c0(w487), .c1(w486), .d0(w1299), .d1(w1300), .x(w1292) );
	dmg_aon2222 g1254 (.a0(w896), .a1(w33), .b0(w32), .b1(w1291), .c0(w889), .c1(w888), .d0(w893), .d1(w894), .x(w41) );
	dmg_notif1 g1255 (.ena(w582), .a(w572), .x(w180) );
	dmg_notif1 g1256 (.ena(w582), .a(w756), .x(w187) );
	dmg_notif1 g1257 (.ena(w582), .a(w757), .x(w229) );
	dmg_notif1 g1258 (.ena(w582), .a(w1155), .x(w29) );
	dmg_notif1 g1259 (.ena(w582), .a(w1156), .x(w16) );
	dmg_notif1 g1260 (.ena(w582), .a(w377), .x(w331) );
	dmg_notif1 g1261 (.ena(w582), .a(w513), .x(w183) );
	dmg_notif1 g1262 (.ena(w582), .a(w645), .x(w55) );
	dmg_not g1263 (.a(w144), .x(w773) );
	dmg_notif0 g1264 (.n_ena(w116), .a(w436), .x(w331) );
	dmg_nand5 g1265 (.a(w134), .b(w133), .c(w129), .d(w1061), .e(w834), .x(w833) );
	dmg_nand5 g1266 (.a(w956), .b(w578), .c(w112), .d(w800), .e(w801), .x(w1199) );
	dmg_nand5 g1267 (.a(w502), .b(w353), .c(w91), .d(w355), .e(w1209), .x(w92) );
	dmg_nand5 g1268 (.a(w439), .b(w440), .c(w156), .d(w541), .e(w471), .x(w470) );
	dmg_not g1269 (.a(w180), .x(w547) );
	dmg_not g1270 (.a(w1296), .x(w1295) );
	dmg_const g1271 (.q0(w20) );
	dmg_xor g1272 (.a(w231), .b(w1001), .x(w1132) );
	dmg_xor g1273 (.a(w231), .b(w306), .x(w1002) );
	dmg_xor g1274 (.a(w231), .b(w301), .x(w300) );
	dmg_xor g1275 (.a(w231), .b(w1078), .x(w868) );
	dmg_xor g1276 (.a(w231), .b(w268), .x(w267) );
	dmg_xor g1277 (.a(w231), .b(w793), .x(w863) );
	dmg_xor g1278 (.a(w231), .b(w862), .x(w859) );
	dmg_xor g1279 (.a(w231), .b(w265), .x(w935) );
	dmg_xor g1280 (.a(w231), .b(w794), .x(w266) );
	dmg_xor g1281 (.a(w231), .b(w871), .x(w416) );
	dmg_and3 g1282 (.a(w1082), .b(w1081), .c(w1022), .x(w1023) );
	dmg_and3 g1283 (.a(w288), .b(w290), .c(w289), .x(w308) );
	dmg_and3 g1284 (.a(w941), .b(w309), .c(w1076), .x(w1133) );
	dmg_and3 g1285 (.a(w292), .b(w1310), .c(w1089), .x(w1033) );
	dmg_and3 g1286 (.a(w611), .b(w723), .c(w454), .x(w556) );
	dmg_and3 g1287 (.a(w372), .b(w373), .c(w1234), .x(w1229) );
	dmg_xor g1288 (.a(w231), .b(w232), .x(w875) );
	dmg_and3 g1289 (.a(w605), .b(w732), .c(w676), .x(w677) );
	dmg_and g1290 (.a(w904), .b(w188), .x(w650) );
	dmg_and g1291 (.a(w933), .b(w932), .x(w1350) );
	dmg_and g1292 (.a(w292), .b(w1310), .x(w1088) );
	dmg_not4 g1293 (.a(w140), .x(w141) );
	dmg_and3 g1294 (.a(w1368), .b(w333), .c(w1369), .x(w1375) );
	dmg_xnor g1295 (.x(w1376), .a(w477), .b(w478) );
	dmg_nand3 g1296 (.a(w1090), .b(w1080), .c(w940), .x(w1089) );
	dmg_or4 g1297 (.a(w111), .b(w711), .c(w112), .d(w666), .x(w1197) );
	dmg_or4 g1298 (.a(w710), .b(w578), .c(w112), .d(w666), .x(w665) );
	dmg_or4 g1299 (.a(w780), .b(w781), .c(w778), .d(w777), .x(w879) );
	dmg_nor5 g1300 (.a(w134), .b(w1269), .c(w339), .d(w480), .e(w481), .x(w836) );
	dmg_nor5 g1301 (.a(w134), .b(w133), .c(w129), .d(w1061), .e(w834), .x(w614) );
	dmg_nor5 g1302 (.a(w502), .b(w353), .c(w91), .d(w355), .e(w1209), .x(w1208) );
	dmg_nor5 g1303 (.a(w502), .b(w352), .c(w351), .d(w348), .e(w361), .x(w755) );
	dmg_and4 g1304 (.a(w208), .b(w315), .c(w63), .d(w209), .x(w318) );
	dmg_and4 g1305 (.a(w208), .b(w206), .c(w63), .d(w209), .x(w316) );
	dmg_or3 g1306 (.a(w574), .b(w582), .c(w581), .x(w704) );
	dmg_dffrnq_comp g1307 (.nr2(w40), .nr1(w40), .d(w891), .ck(w39), .cck(w644), .q(w892), .nq(w891) );
	dmg_dffrnq_comp g1308 (.nr2(w40), .nr1(w40), .d(w890), .ck(w891), .cck(w892), .q(w889), .nq(w890) );
	dmg_dffrnq_comp g1309 (.nr2(w626), .nr1(w626), .d(w489), .ck(w490), .cck(w491), .q(w488), .nq(w489) );
	dmg_dffrnq_comp g1310 (.nr2(w626), .nr1(w626), .d(w1298), .ck(w489), .cck(w488), .q(w487), .nq(w1298) );
	dmg_not g1311 (.a(w491), .x(w492) );
	dmg_or3 g1312 (.a(w70), .b(w507), .c(w755), .x(w923) );
	dmg_or3 g1313 (.a(w70), .b(w1195), .c(w408), .x(w407) );
	dmg_or3 g1314 (.a(w679), .b(w681), .c(w682), .x(w673) );
	dmg_or3 g1315 (.a(w369), .b(w428), .c(w427), .x(w434) );
	dmg_or3 g1316 (.a(w809), .b(w977), .c(w978), .x(w135) );
	dmg_or3 g1317 (.a(w70), .b(w1070), .c(w836), .x(w837) );
	dmg_not g1318 (.a(w566), .x(w237) );
	dmg_nor4 g1319 (.a(w856), .b(w977), .c(w340), .d(w70), .x(w341) );
	dmg_nor4 g1320 (.a(w1380), .b(w428), .c(w27), .d(w70), .x(w878) );
	dmg_not g1321 (.a(w369), .x(w368) );
	dmg_nor5 g1322 (.a(w439), .b(w440), .c(w156), .d(w541), .e(w471), .x(w772) );
	dmg_nor5 g1323 (.a(w439), .b(w438), .c(w214), .d(w848), .e(w530), .x(w529) );
	dmg_or g1324 (.a(w822), .b(w44), .x(w483) );
	dmg_nor4 g1325 (.a(w672), .b(w681), .c(w347), .d(w70), .x(w678) );
	dmg_and3 g1326 (.a(w995), .b(w996), .c(w1034), .x(w342) );
	dmg_nor6 g1327 (.a(w666), .b(w111), .c(w110), .d(w104), .e(w103), .f(w667), .x(w1342) );
	dmg_or4 g1328 (.a(w21), .b(w70), .c(w22), .d(w529), .x(w1303) );
	dmg_and4 g1329 (.a(w801), .b(w114), .c(w113), .d(w951), .x(w115) );
endmodule // APU