// 8 bit lanes x 4 cols x 32 rows = 1024 bit

module HRAM (  clk7, soc_rd, soc_wr, d, ffxx, a);

	input wire clk7;
	input wire soc_rd;
	input wire soc_wr;
	inout wire [7:0]d;
	input wire ffxx;
	input wire [7:0]a

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire [31:0]w45;
	wire [3:0]w46;
	wire [3:0]w47;
	wire [3:0]w48;
	wire [3:0]w49;
	wire [3:0]w50;
	wire [3:0]w51;
	wire [3:0]w52;
	wire [3:0]w53;
	wire [3:0]w54;
	wire [3:0]w55;
	wire [3:0]w56;
	wire [3:0]w57;
	wire [3:0]w58;
	wire [3:0]w59;
	wire [3:0]w60;
	wire [3:0]w61;

	assign w34 = clk7;
	assign w35 = soc_rd;
	assign w36 = soc_wr;
	assign d[0] = w37;
	assign d[1] = w38;
	assign d[2] = w39;
	assign d[3] = w40;
	assign d[4] = w41;
	assign d[5] = w42;
	assign d[6] = w43;
	assign d[7] = w44;
	assign w14 = ffxx;
	assign w16 = a[0];
	assign w15 = a[1];
	assign w19 = a[2];
	assign w20 = a[3];
	assign w21 = a[4];
	assign w22 = a[5];
	assign w23 = a[6];
	assign w24 = a[7];

	// Instances

	sram_bit_lane g1 (.db(w39), .n_oe(w10), .n_pch(w9), .oe(w6), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w56), .bl(w57) );
	sram_bit_lane g2 (.db(w40), .n_pch(w9), .n_oe(w10), .oe(w6), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w54), .bl(w55) );
	sram_bit_lane g3 (.db(w41), .oe(w6), .n_pch(w9), .n_oe(w10), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w52), .bl(w53) );
	sram_bit_lane g4 (.db(w42), .n_pch(w9), .n_oe(w10), .oe(w6), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w50), .bl(w51) );
	sram_bit_lane g5 (.db(w43), .oe(w6), .n_pch(w9), .n_oe(w10), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w48), .bl(w49) );
	sram_bit_lane g6 (.db(w44), .oe(w6), .n_pch(w9), .n_oe(w10), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w47), .bl(w46) );
	sram_bit_lane g7 (.db(w37), .oe(w6), .n_pch(w9), .n_oe(w10), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w60), .bl(w61) );
	sram_bit_lane g8 (.db(w38), .oe(w6), .n_pch(w9), .n_oe(w10), .wr(w8), .c[3](w30), .c[2](w33), .c[1](w32), .c[0](w31), .n_bl(w58), .bl(w59) );
	sram_array g9 (.n_pch(w9), .n_BL(w60), .BL(w61), .WL(w45) );
	sram_array g10 (.n_pch(w9), .n_BL(w58), .BL(w59), .WL(w45) );
	sram_array g11 (.n_pch(w9), .n_BL(w56), .BL(w57), .WL(w45) );
	sram_array g12 (.n_pch(w9), .n_BL(w54), .BL(w55), .WL(w45) );
	sram_array g13 (.n_pch(w9), .n_BL(w52), .BL(w53), .WL(w45) );
	sram_array g14 (.n_pch(w9), .n_BL(w50), .BL(w51), .WL(w45) );
	sram_array g15 (.n_pch(w9), .n_BL(w48), .BL(w49), .WL(w45) );
	sram_array g16 (.n_pch(w9), .WL(w45), .n_BL(w47), .BL(w46) );
	dmg_not2 g17 (.a(w7), .x(w9) );
	dmg_not g18 (.a(w6), .x(w10) );
	dmg_not2 g19 (.a(w5), .x(w6) );
	dmg_not2 g20 (.a(w13), .x(w8) );
	dmg_not g21 (.a(w16), .x(w17) );
	dmg_not g22 (.a(w15), .x(w18) );
	dmg_not2 g23 (.a(w1), .x(w11) );
	dmg_not2 g24 (.a(w3), .x(w12) );
	dmg_not g25 (.a(w23), .x(w25) );
	dmg_not g26 (.a(w22), .x(w26) );
	dmg_not g27 (.a(w21), .x(w27) );
	dmg_not g28 (.a(w20), .x(w28) );
	dmg_not g29 (.a(w19), .x(w29) );
	dmg_nand g30 (.b(w9), .a(w2), .x(w1) );
	dmg_or g31 (.b(w8), .a(w6), .x(w2) );
	dmg_nand3 g32 (.c(w14), .b(w24), .a(w4), .x(w3) );
	dmg_nand7 g33 (.g(w23), .f(w22), .e(w21), .d(w20), .c(w19), .b(w15), .a(w16), .x(w4) );
	dmg_and g34 (.a(w16), .b(w15), .x(w30) );
	dmg_and g35 (.a(w17), .b(w15), .x(w33) );
	dmg_and g36 (.a(w18), .b(w16), .x(w32) );
	dmg_and g37 (.a(w17), .b(w18), .x(w31) );
	dmg_nand g38 (.a(w12), .b(w36), .x(w13) );
	dmg_nand g39 (.a(w12), .b(w35), .x(w5) );
	dmg_nor3 g40 (.a(w34), .b(w8), .c(w6), .x(w7) );
	sram_row_decode g41 (.n_wl_pch(w11), .wl_ena(w12), .d[0](w19), .d[1](w20), .d[2](w21), .d[3](w22), .d[4](w23), .nd[0](w29), .nd[1](w28), .nd[2](w27), .nd[3](w26), .nd[4](w25), .x(w45) );
endmodule // HRAM