module APU (  cclk, clk2, clk4, clk6, clk7, clk9, n_reset2, a, d, cpu_wakeup, n_DRV_HIGH_a, n_INPUT_a, DRV_LOW_a,  
	n_sout_topad, n_DRV_HIGH_sin, n_ENA_PU_sin, DRV_LOW_sin, n_DRV_HIGH_sck, sck_dir, DRV_LOW_sck, n_DRV_HIGH_p10, CONST0, n_p10, DRV_LOW_p10, n_DRV_HIGH_p11, n_p11, DRV_LOW_p11, n_DRV_HIGH_p12, n_p12, DRV_LOW_p12, n_DRV_HIGH_p13, n_p13, DRV_LOW_p13, n_DRV_HIGH_p14, DRV_LOW_p14, n_DRV_HIGH_p15, DRV_LOW_p15, 
	dma_a, soc_wr, soc_rd, lfo_512Hz, ser_out, serial_tick, test_1, test_2, n_ext_addr_en, ch3_active, 
	wave_a, wave_rd, n_wave_wr, wave_bl_pch, n_wave_rd, addr_latch, int_jp, FF60_D1, ffxx, n_ch1_amp_en, n_ch2_amp_en, n_ch3_amp_en, n_ch4_amp_en, 
	ch1_out, ch2_out, ch3_out, ch4_out, r_vin_en, rmixer, l_vin_en, lmixer, n_rvolume, n_lvolume, dma_addr_ext);

	input wire cclk;
	input wire clk2;
	input wire clk4;
	input wire clk6;
	input wire clk7;
	input wire clk9;
	input wire n_reset2;
	inout wire [7:0] a; 			// 7:0 are used only   ⚠️ bidir
	inout wire [7:0] d;
	output wire cpu_wakeup;
	output wire [7:0] n_DRV_HIGH_a;
	input wire [7:0] n_INPUT_a;
	output wire [7:0] DRV_LOW_a;
	output wire n_sout_topad;
	output wire n_DRV_HIGH_sin;
	output wire n_ENA_PU_sin;
	output wire DRV_LOW_sin;
	output wire n_DRV_HIGH_sck;
	input wire sck_dir;
	output wire DRV_LOW_sck;
	output wire n_DRV_HIGH_p10;
	inout wire CONST0;
	input wire n_p10;
	output wire DRV_LOW_p10;
	output wire n_DRV_HIGH_p11;
	input wire n_p11;
	output wire DRV_LOW_p11;
	output wire n_DRV_HIGH_p12;
	input wire n_p12;
	output wire DRV_LOW_p12;
	output wire n_DRV_HIGH_p13;
	input wire n_p13;
	output wire DRV_LOW_p13;
	output wire n_DRV_HIGH_p14;
	output wire DRV_LOW_p14;
	output wire n_DRV_HIGH_p15;
	output wire DRV_LOW_p15;
	input wire [7:0] dma_a; 		// 7:0 are used only
	input wire soc_wr;
	input wire soc_rd;
	input wire lfo_512Hz;
	input wire ser_out;
	input wire serial_tick;
	input wire test_1;
	input wire test_2;
	input wire n_ext_addr_en;
	output wire ch3_active;
	output wire [3:0] wave_a;
	input wire [7:0] wave_rd;
	output wire n_wave_wr;
	output wire wave_bl_pch;
	output wire n_wave_rd;
	input wire addr_latch;
	output wire int_jp;
	output wire FF60_D1;
	input wire ffxx;
	output wire n_ch1_amp_en;
	output wire n_ch2_amp_en;
	output wire n_ch3_amp_en;
	output wire n_ch4_amp_en;
	output wire [3:0] ch1_out;
	output wire [3:0] ch2_out;
	output wire [3:0] ch3_out;
	output wire [3:0] ch4_out;
	output wire r_vin_en;
	output wire [3:0] rmixer;
	output wire l_vin_en;
	output wire [3:0] lmixer;
	output wire [2:0] n_rvolume;
	output wire [2:0] n_lvolume;
	input wire dma_addr_ext;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;
	wire w981;
	wire w982;
	wire w983;
	wire w984;
	wire w985;
	wire w986;
	wire w987;
	wire w988;
	wire w989;
	wire w990;
	wire w991;
	wire w992;
	wire w993;
	wire w994;
	wire w995;
	wire w996;
	wire w997;
	wire w998;
	wire w999;
	wire w1000;
	wire w1001;
	wire w1002;
	wire w1003;
	wire w1004;
	wire w1005;
	wire w1006;
	wire w1007;
	wire w1008;
	wire w1009;
	wire w1010;
	wire w1011;
	wire w1012;
	wire w1013;
	wire w1014;
	wire w1015;
	wire w1016;
	wire w1017;
	wire w1018;
	wire w1019;
	wire w1020;
	wire w1021;
	wire w1022;
	wire w1023;
	wire w1024;
	wire w1025;
	wire w1026;
	wire w1027;
	wire w1028;
	wire w1029;
	wire w1030;
	wire w1031;
	wire w1032;
	wire w1033;
	wire w1034;
	wire w1035;
	wire w1036;
	wire w1037;
	wire w1038;
	wire w1039;
	wire w1040;
	wire w1041;
	wire w1042;
	wire w1043;
	wire w1044;
	wire w1045;
	wire w1046;
	wire w1047;
	wire w1048;
	wire w1049;
	wire w1050;
	wire w1051;
	wire w1052;
	wire w1053;
	wire w1054;
	wire w1055;
	wire w1056;
	wire w1057;
	wire w1058;
	wire w1059;
	wire w1060;
	wire w1061;
	wire w1062;
	wire w1063;
	wire w1064;
	wire w1065;
	wire w1066;
	wire w1067;
	wire w1068;
	wire w1069;
	wire w1070;
	wire w1071;
	wire w1072;
	wire w1073;
	wire w1074;
	wire w1075;
	wire w1076;
	wire w1077;
	wire w1078;
	wire w1079;
	wire w1080;
	wire w1081;
	wire w1082;
	wire w1083;
	wire w1084;
	wire w1085;
	wire w1086;
	wire w1087;
	wire w1088;
	wire w1089;
	wire w1090;
	wire w1091;
	wire w1092;
	wire w1093;
	wire w1094;
	wire w1095;
	wire w1096;
	wire w1097;
	wire w1098;
	wire w1099;
	wire w1100;
	wire w1101;
	wire w1102;
	wire w1103;
	wire w1104;
	wire w1105;
	wire w1106;
	wire w1107;
	wire w1108;
	wire w1109;
	wire w1110;
	wire w1111;
	wire w1112;
	wire w1113;
	wire w1114;
	wire w1115;
	wire w1116;
	wire w1117;
	wire w1118;
	wire w1119;
	wire w1120;
	wire w1121;
	wire w1122;
	wire w1123;
	wire w1124;
	wire w1125;
	wire w1126;
	wire w1127;
	wire w1128;
	wire w1129;
	wire w1130;
	wire w1131;
	wire w1132;
	wire w1133;
	wire w1134;
	wire w1135;
	wire w1136;
	wire w1137;
	wire w1138;
	wire w1139;
	wire w1140;
	wire w1141;
	wire w1142;
	wire w1143;
	wire w1144;
	wire w1145;
	wire w1146;
	wire w1147;
	wire w1148;
	wire w1149;
	wire w1150;
	wire w1151;
	wire w1152;
	wire w1153;
	wire w1154;
	wire w1155;
	wire w1156;
	wire w1157;
	wire w1158;
	wire w1159;
	wire w1160;
	wire w1161;
	wire w1162;
	wire w1163;
	wire w1164;
	wire w1165;
	wire w1166;
	wire w1167;
	wire w1168;
	wire w1169;
	wire w1170;
	wire w1171;
	wire w1172;
	wire w1173;
	wire w1174;
	wire w1175;
	wire w1176;
	wire w1177;
	wire w1178;
	wire w1179;
	wire w1180;
	wire w1181;
	wire w1182;
	wire w1183;
	wire w1184;
	wire w1185;
	wire w1186;
	wire w1187;
	wire w1188;
	wire w1189;
	wire w1190;
	wire w1191;
	wire w1192;
	wire w1193;
	wire w1194;
	wire w1195;
	wire w1196;
	wire w1197;
	wire w1198;
	wire w1199;
	wire w1200;
	wire w1201;
	wire w1202;
	wire w1203;
	wire w1204;
	wire w1205;
	wire w1206;
	wire w1207;
	wire w1208;
	wire w1209;
	wire w1210;
	wire w1211;
	wire w1212;
	wire w1213;
	wire w1214;
	wire w1215;
	wire w1216;
	wire w1217;
	wire w1218;
	wire w1219;
	wire w1220;
	wire w1221;
	wire w1222;
	wire w1223;
	wire w1224;
	wire w1225;
	wire w1226;
	wire w1227;
	wire w1228;
	wire w1229;
	wire w1230;
	wire w1231;
	wire w1232;
	wire w1233;
	wire w1234;
	wire w1235;
	wire w1236;
	wire w1237;
	wire w1238;
	wire w1239;
	wire w1240;
	wire w1241;
	wire w1242;
	wire w1243;
	wire w1244;
	wire w1245;
	wire w1246;
	wire w1247;
	wire w1248;
	wire w1249;
	wire w1250;
	wire w1251;
	wire w1252;
	wire w1253;
	wire w1254;
	wire w1255;
	wire w1256;
	wire w1257;
	wire w1258;
	wire w1259;
	wire w1260;
	wire w1261;
	wire w1262;
	wire w1263;
	wire w1264;
	wire w1265;
	wire w1266;
	wire w1267;
	wire w1268;
	wire w1269;
	wire w1270;
	wire w1271;
	wire w1272;
	wire w1273;
	wire w1274;
	wire w1275;
	wire w1276;
	wire w1277;
	wire w1278;
	wire w1279;
	wire w1280;
	wire w1281;
	wire w1282;
	wire w1283;
	wire w1284;
	wire w1285;
	wire w1286;
	wire w1287;
	wire w1288;
	wire w1289;
	wire w1290;
	wire w1291;
	wire w1292;
	wire w1293;
	wire w1294;
	wire w1295;
	wire w1296;
	wire w1297;
	wire w1298;
	wire w1299;
	wire w1300;
	wire w1301;
	wire w1302;
	wire w1303;
	wire w1304;
	wire w1305;
	wire w1306;
	wire w1307;
	wire w1308;
	wire w1309;
	wire w1310;
	wire w1311;
	wire w1312;
	wire w1313;
	wire w1314;
	wire w1315;
	wire w1316;
	wire w1317;
	wire w1318;
	wire w1319;
	wire w1320;
	wire w1321;
	wire w1322;
	wire w1323;
	wire w1324;
	wire w1325;
	wire w1326;
	wire w1327;
	wire w1328;
	wire w1329;
	wire w1330;
	wire w1331;
	wire w1332;
	wire w1333;
	wire w1334;
	wire w1335;
	wire w1336;
	wire w1337;
	wire w1338;
	wire w1339;
	wire w1340;
	wire w1341;
	wire w1342;
	wire w1343;
	wire w1344;
	wire w1345;
	wire w1346;
	wire w1347;
	wire w1348;
	wire w1349;
	wire w1350;
	wire w1351;
	wire w1352;
	wire w1353;
	wire w1354;
	wire w1355;
	wire w1356;
	wire w1357;
	wire w1358;
	wire w1359;
	wire w1360;
	wire w1361;
	wire w1362;
	wire w1363;
	wire w1364;
	wire w1365;
	wire w1366;
	wire w1367;
	wire w1368;
	wire w1369;
	wire w1370;
	wire w1371;
	wire w1372;
	wire w1373;
	wire w1374;
	wire w1375;
	wire w1376;
	wire w1377;
	wire w1378;
	wire w1379;
	wire w1380;
	wire w1381;
	wire w1382;
	wire w1383;
	wire w1384;
	wire w1385;
	wire w1386;
	wire w1387;
	wire w1388;
	wire w1389;
	wire w1390;
	wire w1391;
	wire w1392;
	wire w1393;
	wire w1394;
	wire w1395;
	wire w1396;
	wire w1397;
	wire w1398;
	wire w1399;
	wire w1400;
	wire w1401;
	wire w1402;
	wire w1403;
	wire w1404;
	wire w1405;
	wire w1406;
	wire w1407;

	assign w1156 = n_INPUT_a[5];
	assign n_DRV_HIGH_a[5] = w1157;
	assign DRV_LOW_a[6] = w1258;
	assign DRV_LOW_a[5] = w2;
	assign w1 = n_INPUT_a[4];
	assign w88 = n_INPUT_a[6];
	assign n_DRV_HIGH_a[6] = w1257;
	assign DRV_LOW_a[7] = w89;
	assign w708 = n_INPUT_a[7];
	assign n_DRV_HIGH_a[4] = w709;
	assign DRV_LOW_a[1] = w627;
	assign DRV_LOW_a[4] = w628;
	assign n_DRV_HIGH_a[3] = w1263;
	assign n_DRV_HIGH_a[7] = w1160;
	assign w1159 = n_INPUT_a[3];
	assign DRV_LOW_a[3] = w667;
	assign n_DRV_HIGH_a[2] = w1048;
	assign w666 = n_INPUT_a[2];
	assign DRV_LOW_a[2] = w1049;
	assign n_DRV_HIGH_a[1] = w707;
	assign w706 = n_INPUT_a[1];
	assign w447 = n_INPUT_a[0];
	assign n_DRV_HIGH_a[0] = w126;
	assign DRV_LOW_a[0] = w127;
	assign n_sout_topad = w1247;
	assign n_DRV_HIGH_sin = w811;
	assign DRV_LOW_sin = w809;
	assign n_DRV_HIGH_sck = w889;
	assign DRV_LOW_sck = w1287;
	assign n_ENA_PU_sin = w624;
	assign n_DRV_HIGH_p10 = w945;
	assign DRV_LOW_p10 = w568;
	assign n_DRV_HIGH_p13 = w947;
	assign n_DRV_HIGH_p11 = w884;
	assign DRV_LOW_p13 = w946;
	assign DRV_LOW_p11 = w565;
	assign n_DRV_HIGH_p14 = w566;
	assign DRV_LOW_p14 = w626;
	assign w784 = n_p10;
	assign n_DRV_HIGH_p12 = w438;
	assign w785 = n_p11;
	assign w787 = n_p13;
	assign DRV_LOW_p12 = w883;
	assign w788 = n_p12;
	assign DRV_LOW_p15 = w804;
	assign n_DRV_HIGH_p15 = w839;
	assign n_lvolume[2] = w224;
	assign n_rvolume[2] = w1165;
	assign n_rvolume[1] = w378;
	assign n_lvolume[1] = w1163;
	assign n_rvolume[0] = w227;
	assign n_lvolume[0] = w226;
	assign l_vin_en = w1121;
	assign ch4_out[3] = w1164;
	assign ch4_out[2] = w131;
	assign ch4_out[1] = w130;
	assign lmixer[1] = w1082;
	assign ch4_out[0] = w1081;
	assign lmixer[0] = w1106;
	assign rmixer[1] = w1120;
	assign r_vin_en = w822;
	assign lmixer[2] = w1056;
	assign rmixer[2] = w823;
	assign lmixer[3] = w1057;
	assign rmixer[3] = w17;
	assign rmixer[0] = w18;
	assign n_ch4_amp_en = w843;
	assign CONST0 = w20;
	assign ch2_out[3] = w1358;
	assign ch2_out[2] = w1359;
	assign ch2_out[1] = w1342;
	assign n_ch1_amp_en = w533;
	assign ch2_out[0] = w1357;
	assign ch1_out[1] = w549;
	assign w1331 = lfo_512Hz;
	assign ch1_out[0] = w548;
	assign ch1_out[2] = w547;
	assign ch1_out[3] = w546;
	assign w114 = soc_rd;
	assign d[3] = w229;
	assign d[6] = w55;
	assign d[5] = w16;
	assign d[2] = w180;
	assign d[7] = w187;
	assign d[0] = w183;
	assign w807 = soc_wr;
	assign w7 = dma_a[0];
	assign w887 = ffxx;
	assign w888 = sck_dir;
	assign w1214 = clk6;
	assign d[4] = w29;
	assign d[1] = w333;
	assign w8 = clk7;
	assign ch3_out[3] = w720;
	assign ch3_out[2] = w1046;
	assign ch3_out[1] = w1348;
	assign cpu_wakeup = w1215;
	assign a[7] = w672;
	assign w575 = n_reset2;
	assign n_ch2_amp_en = w761;
	assign ch3_out[0] = w760;
	assign w57 = ser_out;
	assign a[6] = w112;
	assign a[4] = w111;
	assign n_ch3_amp_en = w410;
	assign a[2] = w104;
	assign a[5] = w583;
	assign w584 = dma_a[4];
	assign w697 = dma_a[2];
	assign a[3] = w110;
	assign w1344 = test_2;
	assign w11 = clk2;
	assign w10 = clk9;
	assign a[1] = w103;
	assign int_jp = w1047;
	assign w385 = dma_addr_ext;
	assign FF60_D1 = w718;
	assign w387 = dma_a[7];
	assign w388 = cclk;
	assign a[0] = w673;
	assign w1138 = serial_tick;
	assign w1137 = dma_a[3];
	assign w1355 = dma_a[5];
	assign w581 = dma_a[6];
	assign w383 = dma_a[1];
	assign w382 = wave_rd[4];
	assign n_wave_wr = w580;
	assign w1169 = wave_rd[5];
	assign w5 = addr_latch;
	assign n_wave_rd = w711;
	assign w589 = wave_rd[7];
	assign w590 = wave_rd[3];
	assign w405 = wave_rd[1];
	assign wave_bl_pch = w1175;
	assign w1174 = wave_rd[6];
	assign w578 = wave_rd[2];
	assign w90 = test_1;
	assign w518 = wave_rd[0];
	assign ch3_active = w399;
	assign w125 = n_ext_addr_en;
	assign wave_a[3] = w1155;
	assign wave_a[2] = w1154;
	assign wave_a[1] = w1354;
	assign wave_a[0] = w1153;
	assign w123 = clk4;

	// Instances

	dmg_not g1 (.a(w1), .x(w124) );
	dmg_not g2 (.a(w390), .x(w968) );
	dmg_not g3 (.a(w390), .x(w969) );
	dmg_not g4 (.a(w1156), .x(w1173) );
	dmg_not g5 (.a(w578), .x(w577) );
	dmg_not g6 (.a(w1170), .x(w714) );
	dmg_not g7 (.a(w416), .x(w523) );
	dmg_not g8 (.a(w390), .x(w1177) );
	dmg_not g9 (.a(w416), .x(w702) );
	dmg_not g10 (.a(w589), .x(w762) );
	dmg_not g11 (.a(w590), .x(w763) );
	dmg_not g12 (.a(w1170), .x(w1171) );
	dmg_not g13 (.a(w710), .x(w712) );
	dmg_not g14 (.a(w388), .x(w389) );
	dmg_not g15 (.a(w416), .x(w40) );
	dmg_not g16 (.a(w965), .x(w1208) );
	dmg_not g17 (.a(w111), .x(w716) );
	dmg_not g18 (.a(w672), .x(w1216) );
	dmg_not g19 (.a(w112), .x(w1212) );
	dmg_not g20 (.a(w11), .x(w12) );
	dmg_not g21 (.a(w8), .x(w585) );
	dmg_not g22 (.a(w112), .x(w113) );
	dmg_not g23 (.a(w939), .x(w940) );
	dmg_not g24 (.a(w70), .x(w1091) );
	dmg_not g25 (.a(w70), .x(w1034) );
	dmg_not g26 (.a(w390), .x(w1060) );
	dmg_not g27 (.a(w76), .x(w223) );
	dmg_not g28 (.a(w70), .x(w1118) );
	dmg_not g29 (.a(w69), .x(w1119) );
	dmg_not g30 (.a(w44), .x(w837) );
	dmg_not g31 (.a(w44), .x(w836) );
	dmg_not g32 (.a(w833), .x(w834) );
	dmg_not g33 (.a(w78), .x(w79) );
	dmg_not g34 (.a(w1036), .x(w1037) );
	dmg_not g35 (.a(w1101), .x(w1035) );
	dmg_not g36 (.a(w283), .x(w284) );
	dmg_not g37 (.a(w166), .x(w167) );
	dmg_not g38 (.a(w292), .x(w1330) );
	dmg_not g39 (.a(w144), .x(w300) );
	dmg_not g40 (.a(w144), .x(w938) );
	dmg_not g41 (.a(w44), .x(w1143) );
	dmg_not g42 (.a(w217), .x(w1321) );
	dmg_not g43 (.a(w83), .x(w288) );
	dmg_not g44 (.a(w1005), .x(w1006) );
	dmg_not g45 (.a(w1319), .x(w1318) );
	dmg_not g46 (.a(w1202), .x(w1201) );
	dmg_not g47 (.a(w167), .x(w168) );
	dmg_not g48 (.a(w951), .x(w1000) );
	dmg_not g49 (.a(w70), .x(w954) );
	dmg_not g50 (.a(w1307), .x(w1308) );
	dmg_not g51 (.a(w1014), .x(w1015) );
	dmg_not g52 (.a(w44), .x(w1188) );
	dmg_not g53 (.a(w65), .x(w66) );
	dmg_not g54 (.a(w416), .x(w632) );
	dmg_not g55 (.a(w971), .x(w1316) );
	dmg_not g56 (.a(w497), .x(w1313) );
	dmg_not g57 (.a(w84), .x(w83) );
	dmg_not g58 (.a(w894), .x(w319) );
	dmg_not g59 (.a(w1219), .x(w38) );
	dmg_not g60 (.a(w88), .x(w997) );
	dmg_not g61 (.a(w708), .x(w87) );
	dmg_not g62 (.a(w405), .x(w379) );
	dmg_not g63 (.a(w381), .x(w380) );
	dmg_not g64 (.a(w518), .x(w517) );
	dmg_not g65 (.a(w555), .x(w652) );
	dmg_not g66 (.a(w1174), .x(w651) );
	dmg_not g67 (.a(w416), .x(w1260) );
	dmg_not g68 (.a(w706), .x(w705) );
	dmg_not g69 (.a(w390), .x(w392) );
	dmg_not g70 (.a(w416), .x(w1334) );
	dmg_not g71 (.a(w416), .x(w1333) );
	dmg_not g72 (.a(w390), .x(w391) );
	dmg_not g73 (.a(w750), .x(w751) );
	dmg_not g74 (.a(w1226), .x(w1227) );
	dmg_not g75 (.a(w1255), .x(w1304) );
	dmg_not g76 (.a(w555), .x(w554) );
	dmg_not g77 (.a(w408), .x(w407) );
	dmg_not g78 (.a(w399), .x(w400) );
	dmg_not g79 (.a(w923), .x(w170) );
	dmg_not g80 (.a(w70), .x(w152) );
	dmg_not g81 (.a(w229), .x(w1196) );
	dmg_not g82 (.a(w144), .x(w771) );
	dmg_not g83 (.a(w322), .x(w321) );
	dmg_not g84 (.a(w845), .x(w1381) );
	dmg_not g85 (.a(w42), .x(w43) );
	dmg_not g86 (.a(w828), .x(w1372) );
	dmg_not g87 (.a(w480), .x(w119) );
	dmg_not g88 (.a(w119), .x(w118) );
	dmg_not g89 (.a(w816), .x(w815) );
	dmg_not g90 (.a(w865), .x(w864) );
	dmg_not g91 (.a(w326), .x(w327) );
	dmg_not g92 (.a(w830), .x(w477) );
	dmg_not g93 (.a(w893), .x(w829) );
	dmg_not g94 (.a(w151), .x(w892) );
	dmg_not g95 (.a(w333), .x(w329) );
	dmg_not g96 (.a(w70), .x(w121) );
	dmg_not g97 (.a(w1206), .x(w1205) );
	dmg_not g98 (.a(w70), .x(w1204) );
	dmg_not g99 (.a(w926), .x(w925) );
	dmg_not g100 (.a(w1295), .x(w1294) );
	dmg_not g101 (.a(w923), .x(w924) );
	dmg_not g102 (.a(w541), .x(w542) );
	dmg_not g103 (.a(w923), .x(w1233) );
	dmg_not g104 (.a(w44), .x(w1235) );
	dmg_not g105 (.a(w210), .x(w1234) );
	dmg_not g106 (.a(w44), .x(w504) );
	dmg_not g107 (.a(w1142), .x(w1290) );
	dmg_not g108 (.a(w909), .x(w1267) );
	dmg_not g109 (.a(w44), .x(w402) );
	dmg_not g110 (.a(w508), .x(w727) );
	dmg_not g111 (.a(w505), .x(w1353) );
	dmg_not g112 (.a(w70), .x(w1368) );
	dmg_not g113 (.a(w1369), .x(w1370) );
	dmg_not g114 (.a(w555), .x(w459) );
	dmg_not g115 (.a(w529), .x(w556) );
	dmg_not g116 (.a(w1396), .x(w1397) );
	dmg_not g117 (.a(w560), .x(w559) );
	dmg_not g118 (.a(w685), .x(w686) );
	dmg_not g119 (.a(w604), .x(w744) );
	dmg_not g120 (.a(w70), .x(w600) );
	dmg_not g121 (.a(w70), .x(w606) );
	dmg_not g122 (.a(w1274), .x(w665) );
	dmg_not g123 (.a(w347), .x(w741) );
	dmg_not g124 (.a(w609), .x(w610) );
	dmg_not g125 (.a(w368), .x(w367) );
	dmg_not g126 (.a(w680), .x(w681) );
	dmg_not g127 (.a(w44), .x(w736) );
	dmg_not g128 (.a(w44), .x(w729) );
	dmg_not g129 (.a(w70), .x(w365) );
	dmg_not g130 (.a(w965), .x(w1289) );
	dmg_not g131 (.a(w1237), .x(w1236) );
	dmg_not g132 (.a(w16), .x(w1246) );
	dmg_not g133 (.a(w624), .x(w1245) );
	dmg_not g134 (.a(w888), .x(w1244) );
	dmg_not g135 (.a(w867), .x(w271) );
	dmg_not g136 (.a(w233), .x(w236) );
	dmg_not g137 (.a(w480), .x(w1404) );
	dmg_not g138 (.a(w1019), .x(w1020) );
	dmg_not g139 (.a(w48), .x(w1021) );
	dmg_not g140 (.a(w1021), .x(w1022) );
	dmg_not g141 (.a(w44), .x(w1406) );
	dmg_not g142 (.a(w42), .x(w45) );
	dmg_not g143 (.a(w44), .x(w338) );
	dmg_not g144 (.a(w336), .x(w337) );
	dmg_not g145 (.a(w241), .x(w139) );
	dmg_not g146 (.a(w50), .x(w49) );
	dmg_not g147 (.a(w118), .x(w50) );
	dmg_not g148 (.a(w781), .x(w782) );
	dmg_not g149 (.a(w255), .x(w872) );
	dmg_not g150 (.a(w233), .x(w234) );
	dmg_not g151 (.a(w233), .x(w941) );
	dmg_not g152 (.a(w144), .x(w471) );
	dmg_not g153 (.a(w372), .x(w373) );
	dmg_not g154 (.a(w257), .x(w256) );
	dmg_not g155 (.a(w624), .x(w567) );
	dmg_not g156 (.a(w44), .x(w1349) );
	dmg_not g157 (.a(w1238), .x(w1237) );
	dmg_not g158 (.a(w730), .x(w1241) );
	dmg_not g159 (.a(w70), .x(w1240) );
	dmg_not g160 (.a(w29), .x(w469) );
	dmg_not g161 (.a(w447), .x(w446) );
	dmg_not g162 (.a(w70), .x(w731) );
	dmg_not g163 (.a(w468), .x(w732) );
	dmg_not g164 (.a(w203), .x(w202) );
	dmg_not g165 (.a(w732), .x(w733) );
	dmg_not g166 (.a(w70), .x(w194) );
	dmg_not g167 (.a(w70), .x(w461) );
	dmg_not g168 (.a(w454), .x(w453) );
	dmg_not g169 (.a(w465), .x(w464) );
	dmg_not g170 (.a(w70), .x(w197) );
	dmg_not g171 (.a(w347), .x(w196) );
	dmg_not g172 (.a(w347), .x(w198) );
	dmg_not g173 (.a(w186), .x(w185) );
	dmg_not g174 (.a(w1273), .x(w1274) );
	dmg_not g175 (.a(w608), .x(w607) );
	dmg_not g176 (.a(w181), .x(w182) );
	dmg_not g177 (.a(w70), .x(w755) );
	dmg_not g178 (.a(w455), .x(w913) );
	dmg_not g179 (.a(w70), .x(w433) );
	dmg_not g180 (.a(w965), .x(w966) );
	dmg_not g181 (.a(w70), .x(w1231) );
	dmg_not g182 (.a(w210), .x(w211) );
	dmg_not g183 (.a(w144), .x(w774) );
	dmg_not g184 (.a(w473), .x(w472) );
	dmg_not g185 (.a(w860), .x(w861) );
	dmg_not g186 (.a(w571), .x(w799) );
	dmg_not g187 (.a(w796), .x(w797) );
	dmg_not g188 (.a(w1373), .x(w1374) );
	dmg_not g189 (.a(w70), .x(w52) );
	dmg_not g190 (.a(w136), .x(w137) );
	dmg_not g191 (.a(w70), .x(w340) );
	dmg_not g192 (.a(w322), .x(w72) );
	dmg_not g193 (.a(w44), .x(w827) );
	dmg_not g194 (.a(w70), .x(w263) );
	dmg_not g195 (.a(w219), .x(w218) );
	dmg_not g196 (.a(w881), .x(w880) );
	dmg_not g197 (.a(w161), .x(w852) );
	dmg_not g198 (.a(w411), .x(w412) );
	dmg_not g199 (.a(w1292), .x(w1291) );
	dmg_not g200 (.a(w70), .x(w513) );
	dmg_not g201 (.a(w909), .x(w908) );
	dmg_not g202 (.a(w92), .x(w93) );
	dmg_not g203 (.a(w911), .x(w912) );
	dmg_not g204 (.a(w1265), .x(w552) );
	dmg_not g205 (.a(w180), .x(w531) );
	dmg_not g206 (.a(w644), .x(w1264) );
	dmg_not g207 (.a(w692), .x(w1302) );
	dmg_not g208 (.a(w1275), .x(w690) );
	dmg_not g209 (.a(w665), .x(w752) );
	dmg_not g210 (.a(w100), .x(w101) );
	dmg_not g211 (.a(w407), .x(w406) );
	dmg_not g212 (.a(w1184), .x(w1162) );
	dmg_not g213 (.a(w1304), .x(w1219) );
	dmg_not g214 (.a(w44), .x(w1132) );
	dmg_not g215 (.a(w650), .x(w902) );
	dmg_not g216 (.a(w32), .x(w900) );
	dmg_not g217 (.a(w55), .x(w31) );
	dmg_not g218 (.a(w630), .x(w631) );
	dmg_not g219 (.a(w183), .x(w516) );
	dmg_not g220 (.a(w1187), .x(w1186) );
	dmg_not g221 (.a(w168), .x(w169) );
	dmg_not g222 (.a(w514), .x(w515) );
	dmg_not g223 (.a(w70), .x(w972) );
	dmg_not g224 (.a(w932), .x(w973) );
	dmg_not g225 (.a(w187), .x(w769) );
	dmg_not g226 (.a(w770), .x(w974) );
	dmg_not g227 (.a(w1191), .x(w1192) );
	dmg_not g228 (.a(w161), .x(w160) );
	dmg_not g229 (.a(w919), .x(w917) );
	dmg_not g230 (.a(w161), .x(w920) );
	dmg_not g231 (.a(w322), .x(w323) );
	dmg_not g232 (.a(w977), .x(w976) );
	dmg_not g233 (.a(w287), .x(w286) );
	dmg_not g234 (.a(w219), .x(w281) );
	dmg_not g235 (.a(w840), .x(w621) );
	dmg_not g236 (.a(w846), .x(w845) );
	dmg_not g237 (.a(w994), .x(w995) );
	dmg_not g238 (.a(w70), .x(w1055) );
	dmg_not g239 (.a(w44), .x(w1103) );
	dmg_not g240 (.a(w298), .x(w1053) );
	dmg_not g241 (.a(w314), .x(w313) );
	dmg_not g242 (.a(w1324), .x(w21) );
	dmg_not g243 (.a(w333), .x(w1361) );
	dmg_not g244 (.a(w183), .x(w1362) );
	dmg_not g245 (.a(w283), .x(w282) );
	dmg_not g246 (.a(w115), .x(w116) );
	dmg_not g247 (.a(w44), .x(w1110) );
	dmg_not g248 (.a(w1044), .x(w1109) );
	dmg_not g249 (.a(w893), .x(w1111) );
	dmg_not g250 (.a(w952), .x(w953) );
	dmg_not g251 (.a(w583), .x(w959) );
	dmg_not g252 (.a(w807), .x(w806) );
	dmg_not g253 (.a(w887), .x(w1210) );
	dmg_not g254 (.a(w956), .x(w955) );
	dmg_not g255 (.a(w956), .x(w960) );
	dmg_not g256 (.a(w957), .x(w958) );
	dmg_not g257 (.a(w956), .x(w1278) );
	dmg_not g258 (.a(w1217), .x(w957) );
	dmg_not g259 (.a(w416), .x(w59) );
	dmg_not g260 (.a(w44), .x(w414) );
	dmg_not g261 (.a(w583), .x(w717) );
	dmg_not g262 (.a(w1134), .x(w669) );
	dmg_not g263 (.a(w44), .x(w1133) );
	dmg_not g264 (.a(w1169), .x(w1168) );
	dmg_not g265 (.a(w382), .x(w1167) );
	dmg_not g266 (.a(w1170), .x(w576) );
	dmg_not g267 (.a(w764), .x(w1347) );
	dmg_not g268 (.a(w381), .x(w759) );
	dmg_not g269 (.a(w381), .x(w520) );
	dmg_not g270 (.a(w381), .x(w519) );
	dmg_not g271 (.a(w97), .x(w98) );
	dmg_not g272 (.a(w416), .x(w703) );
	dmg_not g273 (.a(w1159), .x(w695) );
	dmg_not g274 (.a(w666), .x(w1158) );
	dmg_not g275 (.a(w416), .x(w694) );
	dmg_not g276 (.a(w416), .x(w1147) );
	dmg_not g277 (.a(w1149), .x(w1150) );
	dmg_not g278 (.a(w416), .x(w1152) );
	dmg_dffr g279 (.clk(w968), .nr1(w1147), .nr2(w1147), .d(w1148), .q(w1149), .nq(w1148) );
	dmg_dffr g280 (.clk(w969), .nr1(w703), .nr2(w703), .d(w395), .q(w396) );
	dmg_dffr g281 (.clk(w390), .nr2(w703), .d(w394), .q(w395), .nq(w704), .nr1(w703) );
	dmg_dffr g282 (.clk(w1177), .nr1(w702), .nr2(w702), .d(w1178), .q(w283), .nq(w1178) );
	dmg_dffr g283 (.clk(w1208), .nr1(w59), .nr2(w59), .d(w58), .q(w1217), .nq(w58) );
	dmg_dffr g284 (.clk(w1211), .nr1(w575), .nr2(w575), .d(w333), .q(w718) );
	dmg_dffr g285 (.clk(w10), .nr1(w575), .nr2(w575), .d(w9), .q(w719) );
	dmg_dffr g286 (.clk(w10), .nr1(w575), .nr2(w575), .d(w963), .q(w9) );
	dmg_dffr g287 (.clk(w10), .nr1(w575), .nr2(w575), .d(w805), .q(w963) );
	dmg_dffr g288 (.clk(w1060), .nr1(w1055), .nr2(w1055), .d(w1059), .nq(w1059) );
	dmg_dffr g289 (.clk(w1059), .nr1(w1055), .nr2(w1055), .d(w1107), .q(w846), .nq(w1107) );
	dmg_dffr g290 (.clk(w994), .nr1(w825), .nr2(w825), .d(w1124), .q(w1027), .nq(w1124) );
	dmg_dffr g291 (.clk(w285), .nr1(w1034), .nr2(w1034), .d(w1033), .nq(w1033) );
	dmg_dffr g292 (.clk(w1201), .nr1(w164), .nr2(w164), .d(w165), .q(w166), .nq(w165) );
	dmg_dffr g293 (.clk(w574), .nr1(w575), .nr2(w575), .d(w16), .nq(w804) );
	dmg_dffr g294 (.clk(w282), .nr1(w950), .nr2(w950), .d(w296), .nq(w296) );
	dmg_dffr g295 (.clk(w1279), .nr1(w26), .nr2(w26), .d(w25), .q(w24), .nq(w25) );
	dmg_dffr g296 (.clk(w38), .nr1(w40), .nr2(w40), .d(w39), .q(w650), .nq(w39) );
	dmg_dffr g297 (.clk(w1179), .nr1(w1181), .nr2(w1181), .d(w1180), .q(w766), .nq(w1180) );
	dmg_dffr g298 (.clk(w1256), .nr1(w1334), .nr2(w1334), .d(w96), .q(w97) );
	dmg_dffr g299 (.clk(w391), .nr1(w694), .nr2(w694), .d(w693), .q(w692), .nq(w693) );
	dmg_dffr g300 (.clk(w1150), .nr1(w1152), .nr2(w1152), .d(w1151), .q(w1256), .nq(w1151) );
	dmg_dffr g301 (.clk(w1256), .nr1(w750), .nr2(w750), .d(w749), .q(w349) );
	dmg_dffr g302 (.clk(w752), .nr1(w108), .nr2(w108), .d(w1276), .q(w525), .nq(w1276) );
	dmg_dffr g303 (.clk(w1276), .nr1(w108), .nr2(w108), .d(w675), .q(w674), .nq(w675) );
	dmg_dffr g304 (.clk(w675), .nr1(w108), .nr2(w108), .d(w107), .q(w102), .nq(w107) );
	dmg_dffr g305 (.clk(w107), .nr1(w108), .nr2(w108), .d(w106), .q(w105), .nq(w106) );
	dmg_dffr g306 (.clk(w106), .nr1(w108), .nr2(w108), .d(w660), .q(w109), .nq(w660) );
	dmg_dffr g307 (.clk(w169), .nr1(w632), .nr2(w632), .d(w494), .q(w495), .nq(w494) );
	dmg_dffr g308 (.clk(w122), .nr1(w972), .nr2(w972), .d(w930), .q(w928) );
	dmg_dffr g309 (.clk(w149), .nr1(w825), .nr2(w825), .d(w851), .q(w850), .nq(w851) );
	dmg_dffr g310 (.clk(w279), .nr1(w825), .nr2(w825), .d(w280), .q(w1017), .nq(w280) );
	dmg_dffr g311 (.clk(w1068), .nr1(w825), .nr2(w825), .d(w1069), .q(w993), .nq(w1069) );
	dmg_dffr g312 (.clk(w1069), .nr1(w1065), .nr2(w1065), .d(w1064), .q(w1063), .nq(w1064) );
	dmg_dffr g313 (.clk(w1381), .nr1(w483), .nr2(w483), .d(w1389), .q(w272) );
	dmg_dffr g314 (.clk(w141), .nr1(w263), .nr2(w263), .d(w71), .q(w1373) );
	dmg_dffr g315 (.clk(w141), .nr1(w263), .nr2(w263), .d(w342), .q(w71) );
	dmg_dffr g316 (.clk(w141), .nr1(w860), .nr2(w860), .d(w862), .q(w342) );
	dmg_dffr g317 (.clk(w122), .nr1(w121), .nr2(w121), .d(w261), .q(w120) );
	dmg_dffr g318 (.clk(w1397), .nr1(w677), .nr2(w677), .d(w1367), .q(w1255), .nq(w1367) );
	dmg_dffr g319 (.clk(w1302), .nr1(w604), .nr2(w604), .d(w743), .q(w348) );
	dmg_dffr g320 (.clk(w1302), .nr1(w606), .nr2(w606), .d(w348), .q(w605) );
	dmg_dffr g321 (.clk(w692), .nr1(w606), .nr2(w606), .d(w605), .q(w1275) );
	dmg_dffr g322 (.clk(w369), .nr1(w684), .nr2(w684), .d(w683), .q(w685) );
	dmg_dffr g323 (.clk(w966), .nr1(w731), .nr2(w731), .d(w1250), .q(w468), .nq(w1250) );
	dmg_dffr g324 (.clk(w574), .nr1(w563), .nr2(w563), .d(w183), .q(w853) );
	dmg_dffr g325 (.clk(w574), .nr1(w563), .nr2(w563), .d(w180), .q(w625) );
	dmg_dffr g326 (.clk(w118), .nr1(w243), .nr2(w243), .d(w250), .q(w248) );
	dmg_dffr g327 (.clk(w118), .nr1(w243), .nr2(w243), .d(w247), .q(w250) );
	dmg_dffr g328 (.clk(w118), .nr1(w243), .nr2(w243), .d(w1380), .q(w791) );
	dmg_dffr g329 (.clk(w118), .nr1(w243), .nr2(w243), .d(w1378), .q(w1379) );
	dmg_dffr g330 (.clk(w845), .nr1(w139), .nr2(w139), .d(w140), .q(w1377), .nq(w140) );
	dmg_dffr g331 (.clk(w1404), .nr1(w243), .nr2(w243), .d(w1390), .q(w51) );
	dmg_dffr g332 (.clk(w49), .nr1(w243), .nr2(w243), .d(w51), .q(w244) );
	dmg_dffr g333 (.clk(w49), .nr1(w243), .nr2(w243), .d(w244), .q(w246) );
	dmg_dffr g334 (.clk(w49), .nr1(w243), .nr2(w243), .d(w246), .q(w245) );
	dmg_dffr g335 (.clk(w49), .nr1(w243), .nr2(w243), .d(w245), .q(w242) );
	dmg_dffr g336 (.clk(w49), .nr1(w243), .nr2(w243), .d(w242), .q(w1378) );
	dmg_dffr g337 (.clk(w371), .nr1(w428), .nr2(w428), .d(w427), .q(w569) );
	dmg_dffr g338 (.clk(w369), .nr1(w885), .nr2(w885), .d(w1243), .q(w371) );
	dmg_dffr g339 (.clk(w574), .nr1(w563), .nr2(w563), .d(w333), .q(w564) );
	dmg_dffr g340 (.clk(w574), .nr1(w563), .nr2(w563), .d(w29), .nq(w626) );
	dmg_dffr g341 (.clk(w574), .nr1(w563), .nr2(w563), .d(w187), .q(w810) );
	dmg_dffr g342 (.clk(w574), .nr1(w563), .nr2(w563), .d(w229), .q(w1395) );
	dmg_dffr g343 (.clk(w574), .nr1(w575), .nr2(w575), .d(w55), .q(w56) );
	dmg_dffr g344 (.clk(w1289), .nr1(w1240), .nr2(w1240), .d(w1239), .q(w1238), .nq(w1239) );
	dmg_dffr g345 (.clk(w607), .nr1(w602), .nr2(w602), .d(w1386), .q(w1273), .nq(w1386) );
	dmg_dffr g346 (.clk(w685), .nr1(w95), .nr2(w95), .d(w94), .q(w739) );
	dmg_dffr g347 (.clk(w1269), .nr1(w1290), .nr2(w1290), .d(w187), .nq(w1249) );
	dmg_dffr g348 (.clk(w118), .nr1(w243), .nr2(w243), .d(w1379), .q(w1380) );
	dmg_dffr g349 (.clk(w480), .nr1(w243), .nr2(w243), .d(w248), .q(w249) );
	dmg_dffr g350 (.clk(w480), .nr1(w243), .nr2(w243), .d(w249), .q(w1392) );
	dmg_dffr g351 (.clk(w480), .nr1(w243), .nr2(w243), .d(w1392), .q(w818) );
	dmg_dffr g352 (.clk(w480), .nr1(w243), .nr2(w243), .d(w818), .q(w481) );
	dmg_dffr g353 (.clk(w480), .nr1(w243), .nr2(w243), .d(w481), .q(w482) );
	dmg_dffr g354 (.clk(w816), .nr1(w1077), .nr2(w1077), .d(w1074), .q(w1281) );
	dmg_dffr g355 (.clk(w826), .nr1(w73), .nr2(w73), .d(w74), .q(w75), .nq(w74) );
	dmg_dffr g356 (.clk(w369), .nr1(w343), .nr2(w343), .d(w344), .q(w816) );
	dmg_dffr g357 (.clk(w162), .nr1(w152), .nr2(w152), .d(w304), .q(w151) );
	dmg_dffr g358 (.clk(w162), .nr1(w152), .nr2(w152), .d(w27), .q(w304) );
	dmg_dffr g359 (.clk(w162), .nr1(w926), .nr2(w926), .d(w927), .q(w27) );
	dmg_dffr g360 (.clk(w498), .nr1(w543), .nr2(w543), .d(w499), .q(w500), .nq(w499) );
	dmg_dffr g361 (.clk(w122), .nr1(w600), .nr2(w600), .d(w599), .q(w601) );
	dmg_dffr g362 (.clk(w660), .nr1(w662), .nr2(w662), .d(w663), .q(w664), .nq(w663) );
	dmg_dffr g363 (.clk(w1256), .nr1(w1334), .nr2(w1334), .d(w349), .q(w96) );
	dmg_dffr g364 (.clk(w122), .nr1(w1333), .nr2(w1333), .d(w1332), .q(w748) );
	dmg_dffr g365 (.clk(w283), .nr1(w1260), .nr2(w1260), .d(w406), .nq(w1259) );
	dmg_dffr g366 (.clk(w1219), .nr1(w40), .nr2(w40), .d(w41), .q(w933) );
	dmg_dffr g367 (.clk(w168), .nr1(w632), .nr2(w632), .d(w1306), .q(w921) );
	dmg_dffr g368 (.clk(w1104), .nr1(w825), .nr2(w825), .d(w149), .q(w220), .nq(w149) );
	dmg_dffr g369 (.clk(w280), .nr1(w825), .nr2(w825), .d(w1104), .q(w278), .nq(w1104) );
	dmg_dffr g370 (.clk(w1029), .nr1(w825), .nr2(w825), .d(w279), .q(w277), .nq(w279) );
	dmg_dffr g371 (.clk(w276), .nr1(w825), .nr2(w825), .d(w1029), .q(w1030), .nq(w1029) );
	dmg_dffr g372 (.clk(w1124), .nr1(w825), .nr2(w825), .d(w1068), .q(w1023), .nq(w1068) );
	dmg_dffr g373 (.clk(w1067), .nr1(w825), .nr2(w825), .d(w276), .q(w275), .nq(w276) );
	dmg_dffr g374 (.clk(w1405), .nr1(w825), .nr2(w825), .d(w1067), .q(w273), .nq(w1067) );
	dmg_dffr g375 (.clk(w1066), .nr1(w825), .nr2(w825), .d(w1405), .q(w848), .nq(w1405) );
	dmg_dffr g376 (.clk(w1064), .nr1(w1065), .nr2(w1065), .d(w1066), .q(w222), .nq(w1066) );
	dmg_dffr g377 (.clk(w284), .nr1(w1034), .nr2(w1034), .d(w1331), .nq(w1095) );
	dmg_dffr g378 (.clk(w1033), .nr1(w1034), .nr2(w1034), .d(w1096), .nq(w1096) );
	dmg_dffr g379 (.clk(w283), .nr1(w1146), .nr2(w1146), .d(w1032), .nq(w143) );
	dmg_dffr g380 (.clk(w283), .nr1(w308), .nr2(w308), .d(w309), .q(w293) );
	dmg_dffr g381 (.clk(w10), .nr1(w575), .nr2(w575), .d(w886), .q(w805) );
	dmg_dffr g382 (.clk(w1211), .nr1(w575), .nr2(w575), .d(w183), .q(w624) );
	dmg_dffr g383 (.clk(w715), .nr1(w19), .nr2(w19), .d(w16), .q(w86) );
	dmg_dffr g384 (.clk(w1178), .nr1(w702), .nr2(w702), .d(w86), .q(w85) );
	dmg_dffr g385 (.clk(w392), .nr1(w703), .nr2(w703), .d(w393), .q(w394) );
	dmg_dffr g386 (.clk(w390), .nr1(w703), .nr2(w703), .d(w665), .q(w393) );
	dmg_cnt g387 (.d(w16), .load(w714), .nq(w1179), .clk(w1172) );
	dmg_cnt g388 (.q(w1031), .d(w948), .load(w1037), .clk(w281) );
	dmg_cnt g389 (.q(w1093), .d(w1092), .load(w1037), .clk(w1031) );
	dmg_cnt g390 (.q(w289), .d(w949), .load(w1330), .clk(w291) );
	dmg_cnt g391 (.q(w291), .d(w310), .load(w1330), .clk(w290) );
	dmg_cnt g392 (.q(w290), .d(w1086), .load(w1330), .clk(w288) );
	dmg_cnt g393 (.d(w229), .load(w323), .nq(w287), .clk(w82) );
	dmg_cnt g394 (.q(w1202), .d(w306), .load(w920), .nq(w832), .clk(w153) );
	dmg_cnt g395 (.q(w1004), .d(w1131), .load(w976), .clk(w1043) );
	dmg_cnt g396 (.q(w1043), .d(w975), .load(w976), .clk(w958) );
	dmg_cnt g397 (.q(w962), .d(w333), .load(w960), .clk(w1343) );
	dmg_cnt g398 (.d(w229), .load(w960), .nq(w971), .clk(w961) );
	dmg_cnt g399 (.q(w1277), .d(w29), .load(w1278), .clk(w1316) );
	dmg_cnt g400 (.q(w1183), .d(w333), .load(w576), .clk(w1182) );
	dmg_cnt g401 (.q(w765), .d(w180), .load(w576), .clk(w1183) );
	dmg_cnt g402 (.d(w229), .load(w576), .nq(w764), .clk(w765) );
	dmg_cnt g403 (.d(w756), .load(w652), .nq(w1226), .clk(w1252) );
	dmg_cnt g404 (.q(w1252), .d(w1253), .load(w652), .nq(w1254), .clk(w659) );
	dmg_cnt g405 (.q(w1182), .d(w183), .load(w576), .clk(w1186) );
	dmg_cnt g406 (.d(w16), .load(w1278), .nq(w1279), .clk(w1277) );
	dmg_cnt g407 (.d(w1005), .load(w160), .nq(w919), .clk(w159) );
	dmg_cnt g408 (.q(w1127), .d(w298), .load(w920), .nq(w918), .clk(w917) );
	dmg_cnt g409 (.q(w153), .d(w939), .load(w920), .nq(w1013), .clk(w1127) );
	dmg_cnt g410 (.d(w16), .load(w321), .nq(w826), .clk(w859) );
	dmg_cnt g411 (.q(w332), .d(w867), .load(w852), .nq(w328), .clk(w327) );
	dmg_cnt g412 (.d(w229), .load(w924), .nq(w1292), .clk(w544) );
	dmg_cnt g413 (.q(w544), .d(w180), .load(w924), .clk(w1387) );
	dmg_cnt g414 (.q(w1293), .d(w183), .load(w924), .clk(w1294) );
	dmg_cnt g415 (.q(w540), .d(w29), .load(w170), .clk(w1291) );
	dmg_cnt g416 (.d(w1371), .load(w554), .nq(w529), .clk(w1352) );
	dmg_cnt g417 (.q(w1350), .d(w1351), .load(w554), .nq(w1335), .clk(w1336) );
	dmg_cnt g418 (.q(w1352), .d(w553), .load(w554), .nq(w745), .clk(w1350) );
	dmg_cnt g419 (.q(w608), .d(w742), .load(w741), .nq(w1272), .clk(w173) );
	dmg_cnt g420 (.q(w611), .d(w639), .load(w367), .clk(w738) );
	dmg_cnt g421 (.q(w738), .d(w366), .load(w367), .clk(w682) );
	dmg_cnt g422 (.q(w682), .d(w735), .load(w367), .clk(w733) );
	dmg_cnt g423 (.q(w1248), .d(w1242), .load(w373), .clk(w1236) );
	dmg_cnt g424 (.q(w538), .d(w255), .load(w160), .nq(w1140), .clk(w256) );
	dmg_cnt g425 (.q(w258), .d(w571), .load(w852), .nq(w573), .clk(w572) );
	dmg_cnt g426 (.q(w1383), .d(w138), .load(w137), .clk(w1022) );
	dmg_cnt g427 (.q(w335), .d(w334), .load(w137), .clk(w1383) );
	dmg_cnt g428 (.q(w1382), .d(w1286), .load(w137), .clk(w335) );
	dmg_cnt g429 (.d(w570), .load(w852), .nq(w257), .clk(w258) );
	dmg_cnt g430 (.q(w375), .d(w1297), .load(w373), .clk(w1248) );
	dmg_cnt g431 (.q(w374), .d(w376), .load(w373), .clk(w375) );
	dmg_cnt g432 (.q(w449), .d(w199), .load(w198), .nq(w178), .clk(w179) );
	dmg_cnt g433 (.q(w179), .d(w451), .load(w198), .nq(w450), .clk(w448) );
	dmg_cnt g434 (.d(w737), .load(w198), .nq(w465), .clk(w449) );
	dmg_cnt g435 (.q(w448), .d(w452), .load(w198), .nq(w640), .clk(w610) );
	dmg_cnt g436 (.q(w641), .d(w467), .load(w196), .nq(w462), .clk(w463) );
	dmg_cnt g437 (.q(w463), .d(w195), .load(w196), .nq(w642), .clk(w466) );
	dmg_cnt g438 (.q(w466), .d(w193), .load(w196), .nq(w192), .clk(w464) );
	dmg_cnt g439 (.d(w377), .load(w196), .clk(w641) );
	dmg_cnt g440 (.q(w1402), .d(w740), .load(w741), .nq(w184), .clk(w185) );
	dmg_cnt g441 (.q(w173), .d(w1300), .load(w741), .nq(w1301), .clk(w1402) );
	dmg_cnt g442 (.q(w1396), .d(w458), .load(w459), .nq(w614), .clk(w613) );
	dmg_cnt g443 (.q(w613), .d(w612), .load(w459), .nq(w1365), .clk(w1366) );
	dmg_cnt g444 (.q(w1366), .d(w460), .load(w459), .nq(w915), .clk(w556) );
	dmg_cnt g445 (.q(w443), .d(w441), .load(w27), .nq(w444), .clk(w445) );
	dmg_cnt g446 (.q(w474), .d(w534), .load(w27), .clk(w854) );
	dmg_cnt g447 (.q(w545), .d(w855), .load(w27), .nq(w537), .clk(w157) );
	dmg_cnt g448 (.q(w158), .d(w881), .load(w160), .nq(w539), .clk(w538) );
	dmg_cnt g449 (.q(w156), .d(w214), .load(w27), .nq(w536), .clk(w535) );
	dmg_cnt g450 (.q(w572), .d(w796), .load(w852), .nq(w331), .clk(w332) );
	dmg_cnt g451 (.q(w1071), .d(w484), .load(w342), .nq(w1282), .clk(w1073) );
	dmg_cnt g452 (.q(w841), .d(w485), .load(w342), .clk(w1072) );
	dmg_cnt g453 (.q(w129), .d(w341), .load(w342), .nq(w1070), .clk(w842) );
	dmg_cnt g454 (.q(w133), .d(w1283), .load(w342), .nq(w988), .clk(w623) );
	dmg_cnt g455 (.q(w859), .d(w29), .load(w321), .clk(w286) );
	dmg_cnt g456 (.q(w81), .d(w333), .load(w323), .clk(w80) );
	dmg_cnt g457 (.q(w159), .d(w770), .load(w160), .nq(w1203), .clk(w158) );
	dmg_cnt g458 (.q(w1387), .d(w333), .load(w924), .clk(w1293) );
	dmg_cnt g459 (.d(w187), .load(w170), .nq(w498), .clk(w171) );
	dmg_cnt g460 (.q(w171), .d(w55), .load(w170), .clk(w1407) );
	dmg_cnt g461 (.q(w1407), .d(w16), .load(w170), .clk(w540) );
	dmg_cnt g462 (.q(w355), .d(w354), .load(w922), .nq(w906), .clk(w907) );
	dmg_cnt g463 (.q(w91), .d(w353), .load(w922), .nq(w904), .clk(w905) );
	dmg_cnt g464 (.q(w357), .d(w350), .load(w349), .nq(w358), .clk(w359) );
	dmg_cnt g465 (.q(w1222), .d(w363), .load(w349), .clk(w364) );
	dmg_cnt g466 (.q(w1336), .d(w1303), .load(w554), .nq(w1337), .clk(w1227) );
	dmg_cnt g467 (.q(w747), .d(w754), .load(w652), .nq(w753), .clk(w101) );
	dmg_cnt g468 (.q(w659), .d(w658), .load(w652), .nq(w746), .clk(w747) );
	dmg_cnt g469 (.q(w1003), .d(w1002), .load(w976), .clk(w1004) );
	dmg_cnt g470 (.q(w82), .d(w180), .load(w323), .clk(w81) );
	dmg_cnt g471 (.q(w80), .d(w183), .load(w323), .clk(w79) );
	dmg_cnt g472 (.q(w1094), .d(w1102), .load(w1037), .clk(w1093) );
	dmg_cnt g473 (.q(w1343), .d(w183), .load(w960), .clk(w1308) );
	dmg_cnt g474 (.q(w961), .d(w180), .load(w960), .clk(w962) );
	dmg_cnt g475 (.q(w1172), .d(w29), .load(w714), .clk(w1347) );
	dmg_latchr_comp g476 (.n_ena(w230), .d(w29), .ena(w142), .nres(w950), .nq(w1086) );
	dmg_latchr_comp g477 (.n_ena(w230), .d(w229), .ena(w142), .nres(w950), .nq(w1090) );
	dmg_latchr_comp g478 (.n_ena(w1089), .d(w180), .ena(w142), .nres(w1091), .nq(w1102) );
	dmg_latchr_comp g479 (.n_ena(w1089), .d(w333), .ena(w142), .nres(w1091), .nq(w1092) );
	dmg_latchr_comp g480 (.n_ena(w1116), .d(w183), .ena(w996), .nres(w19), .q(w18), .nq(w1166) );
	dmg_latchr_comp g481 (.n_ena(w1116), .d(w229), .ena(w996), .nres(w19), .q(w17), .nq(w820) );
	dmg_latchr_comp g482 (.n_ena(w1115), .d(w183), .ena(w228), .nres(w19), .nq(w227) );
	dmg_latchr_comp g483 (.n_ena(w1115), .d(w229), .ena(w228), .nres(w19), .q(w822), .nq(w821) );
	dmg_latchr_comp g484 (.n_ena(w1115), .d(w180), .ena(w228), .nres(w19), .nq(w1165) );
	dmg_latchr_comp g485 (.n_ena(w1084), .d(w55), .ena(w1085), .nres(w19), .nq(w224) );
	dmg_latchr_comp g486 (.n_ena(w69), .d(w55), .ena(w1119), .nres(w1118), .q(w76), .nq(w77) );
	dmg_latchr_comp g487 (.n_ena(w631), .d(w55), .ena(w630), .nres(w632), .q(w489), .nq(w488) );
	dmg_latchr_comp g488 (.n_ena(w759), .d(w405), .ena(w381), .nres(w523), .nq(w757) );
	dmg_latchr_comp g489 (.n_ena(w759), .d(w1169), .ena(w381), .nres(w523), .nq(w758) );
	dmg_latchr_comp g490 (.n_ena(w519), .d(w518), .ena(w381), .nres(w523), .nq(w526) );
	dmg_latchr_comp g491 (.n_ena(w519), .d(w382), .ena(w381), .nres(w523), .nq(w1261) );
	dmg_latchr_comp g492 (.n_ena(w1184), .d(w187), .ena(w1162), .nres(w1398), .q(w1332) );
	dmg_latchr_comp g493 (.n_ena(w514), .d(w55), .ena(w515), .nres(w513), .q(w512), .nq(w510) );
	dmg_latchr_comp g494 (.n_ena(w1192), .d(w333), .ena(w1191), .nres(w340), .q(w1130), .nq(w1131) );
	dmg_latchr_comp g495 (.n_ena(w1192), .d(w180), .ena(w1191), .nres(w340), .q(w1194), .nq(w1002) );
	dmg_latchr_comp g496 (.n_ena(w1192), .d(w183), .ena(w1191), .nres(w340), .q(w1129), .nq(w975) );
	dmg_latchr_comp g497 (.n_ena(w339), .d(w55), .ena(w817), .nres(w340), .q(w484), .nq(w54) );
	dmg_latchr_comp g498 (.n_ena(w339), .d(w16), .ena(w817), .nres(w340), .q(w341), .nq(w1384) );
	dmg_latchr_comp g499 (.n_ena(w339), .d(w187), .ena(w817), .nres(w340), .q(w485), .nq(w486) );
	dmg_latchr_comp g500 (.n_ena(w339), .d(w229), .ena(w817), .nres(w340), .q(w134), .nq(w622) );
	dmg_latchr_comp g501 (.n_ena(w339), .d(w29), .ena(w817), .nres(w340), .q(w1283), .nq(w1284) );
	dmg_latchr_comp g502 (.n_ena(w982), .d(w55), .ena(w983), .nres(w825), .q(w1025), .nq(w1123) );
	dmg_latchr_comp g503 (.n_ena(w982), .d(w187), .ena(w983), .nres(w825), .q(w981), .nq(w479) );
	dmg_latchr_comp g504 (.n_ena(w1205), .d(w187), .ena(w1206), .nres(w1204), .q(w411), .nq(w410) );
	dmg_latchr_comp g505 (.n_ena(w728), .d(w16), .ena(w1225), .nres(w365), .q(w353), .nq(w352) );
	dmg_latchr_comp g506 (.n_ena(w728), .d(w55), .ena(w1225), .nres(w365), .q(w350), .nq(w351) );
	dmg_latchr_comp g507 (.n_ena(w728), .d(w29), .ena(w1225), .nres(w365), .q(w354), .nq(w561) );
	dmg_latchr_comp g508 (.n_ena(w728), .d(w187), .ena(w1225), .nres(w365), .q(w363), .nq(w362) );
	dmg_latchr_comp g509 (.n_ena(w552), .d(w187), .ena(w1265), .nres(w755), .q(w1371) );
	dmg_latchr_comp g510 (.n_ena(w552), .d(w55), .ena(w1265), .nres(w755), .q(w553) );
	dmg_latchr_comp g511 (.n_ena(w552), .d(w16), .ena(w1265), .nres(w755), .q(w1351) );
	dmg_latchr_comp g512 (.n_ena(w557), .d(w187), .ena(w558), .nres(w598), .q(w599) );
	dmg_latchr_comp g513 (.n_ena(w182), .d(w333), .ena(w181), .nres(w197), .q(w1300) );
	dmg_latchr_comp g514 (.n_ena(w182), .d(w183), .ena(w181), .nres(w197), .q(w740) );
	dmg_latchr_comp g515 (.n_ena(w182), .d(w180), .ena(w181), .nres(w197), .q(w742) );
	dmg_latchr_comp g516 (.n_ena(w453), .d(w183), .ena(w454), .nres(w461), .q(w460) );
	dmg_latchr_comp g517 (.n_ena(w453), .d(w180), .ena(w454), .nres(w461), .q(w458) );
	dmg_latchr_comp g518 (.n_ena(w453), .d(w333), .ena(w454), .nres(w461), .q(w612) );
	dmg_latchr_comp g519 (.n_ena(w201), .d(w333), .ena(w200), .nres(w194), .q(w451) );
	dmg_latchr_comp g520 (.n_ena(w201), .d(w29), .ena(w200), .nres(w194), .q(w193) );
	dmg_latchr_comp g521 (.n_ena(w201), .d(w229), .ena(w200), .nres(w194), .q(w737) );
	dmg_latchr_comp g522 (.n_ena(w201), .d(w180), .ena(w200), .nres(w194), .q(w199) );
	dmg_latchr_comp g523 (.n_ena(w202), .d(w16), .ena(w203), .nres(w194), .q(w195) );
	dmg_latchr_comp g524 (.n_ena(w1241), .d(w183), .ena(w730), .nres(w433), .q(w1299), .nq(w1242) );
	dmg_latchr_comp g525 (.n_ena(w1241), .d(w180), .ena(w730), .nres(w433), .q(w432), .nq(w376) );
	dmg_latchr_comp g526 (.n_ena(w1241), .d(w333), .ena(w730), .nres(w433), .q(w1298), .nq(w1297) );
	dmg_latchr_comp g527 (.n_ena(w858), .d(w16), .ena(w1296), .nres(w433), .q(w214), .nq(w213) );
	dmg_latchr_comp g528 (.n_ena(w858), .d(w29), .ena(w1296), .nres(w433), .q(w441), .nq(w857) );
	dmg_latchr_comp g529 (.n_ena(w858), .d(w55), .ena(w1296), .nres(w433), .q(w855), .nq(w856) );
	dmg_latchr_comp g530 (.n_ena(w858), .d(w229), .ena(w1296), .nres(w433), .q(w442), .nq(w436) );
	dmg_latchr_comp g531 (.n_ena(w858), .d(w187), .ena(w1296), .nres(w433), .q(w534), .nq(w434) );
	dmg_latchr_comp g532 (.n_ena(w1391), .d(w333), .ena(w1285), .nres(w139), .nq(w334) );
	dmg_latchr_comp g533 (.n_ena(w1391), .d(w180), .ena(w1285), .nres(w139), .nq(w1286) );
	dmg_latchr_comp g534 (.n_ena(w1391), .d(w183), .ena(w1285), .nres(w139), .nq(w138) );
	dmg_latchr_comp g535 (.n_ena(w336), .d(w229), .ena(w337), .nres(w52), .q(w790), .nq(w789) );
	dmg_latchr_comp g536 (.n_ena(w202), .d(w55), .ena(w203), .nres(w194), .q(w467) );
	dmg_latchr_comp g537 (.n_ena(w202), .d(w187), .ena(w203), .nres(w194), .q(w377) );
	dmg_latchr_comp g538 (.n_ena(w201), .d(w183), .ena(w200), .nres(w194), .q(w452) );
	dmg_latchr_comp g539 (.n_ena(w1370), .d(w16), .ena(w1369), .nres(w1368), .q(w597), .nq(w594) );
	dmg_latchr_comp g540 (.n_ena(w1370), .d(w55), .ena(w1369), .nres(w1368), .q(w595), .nq(w596) );
	dmg_latchr_comp g541 (.n_ena(w681), .d(w333), .ena(w680), .nres(w365), .q(w1271), .nq(w366) );
	dmg_latchr_comp g542 (.n_ena(w681), .d(w180), .ena(w680), .nres(w365), .q(w1270), .nq(w639) );
	dmg_latchr_comp g543 (.n_ena(w681), .d(w183), .ena(w680), .nres(w365), .q(w734), .nq(w735) );
	dmg_latchr_comp g544 (.n_ena(w541), .d(w55), .ena(w542), .nres(w1231), .q(w501), .nq(w502) );
	dmg_latchr_comp g545 (.n_ena(w828), .d(w187), .ena(w1372), .nres(w262), .q(w261) );
	dmg_latchr_comp g546 (.n_ena(w982), .d(w29), .ena(w983), .nres(w825), .q(w990), .nq(w979) );
	dmg_latchr_comp g547 (.n_ena(w982), .d(w16), .ena(w983), .nres(w825), .q(w991), .nq(w980) );
	dmg_latchr_comp g548 (.n_ena(w728), .d(w229), .ena(w1225), .nres(w365), .q(w506), .nq(w360) );
	dmg_latchr_comp g549 (.n_ena(w1264), .d(w1266), .ena(w644), .nres(w19), .q(w1038), .nq(w1223) );
	dmg_latchr_comp g550 (.n_ena(w657), .d(w29), .ena(w656), .nres(w755), .q(w1303) );
	dmg_latchr_comp g551 (.n_ena(w657), .d(w229), .ena(w656), .nres(w755), .q(w756) );
	dmg_latchr_comp g552 (.n_ena(w657), .d(w180), .ena(w656), .nres(w755), .q(w1253) );
	dmg_latchr_comp g553 (.n_ena(w657), .d(w333), .ena(w656), .nres(w755), .q(w658) );
	dmg_latchr_comp g554 (.n_ena(w657), .d(w183), .ena(w656), .nres(w755), .q(w754) );
	dmg_latchr_comp g555 (.n_ena(w631), .d(w187), .ena(w630), .nres(w632), .q(w635), .nq(w636) );
	dmg_latchr_comp g556 (.n_ena(w1014), .d(w187), .ena(w1015), .nres(w929), .q(w930) );
	dmg_latchr_comp g557 (.n_ena(w1115), .d(w333), .ena(w228), .nres(w19), .nq(w378) );
	dmg_latchr_comp g558 (.n_ena(w1116), .d(w333), .ena(w996), .nres(w19), .q(w1120), .nq(w1117) );
	dmg_latchr_comp g559 (.n_ena(w1116), .d(w180), .ena(w996), .nres(w19), .q(w823), .nq(w824) );
	dmg_latchr_comp g560 (.n_ena(w1084), .d(w16), .ena(w1085), .nres(w19), .nq(w1163) );
	dmg_latchr_comp g561 (.n_ena(w1084), .d(w187), .ena(w1085), .nres(w19), .q(w1121), .nq(w1122) );
	dmg_latchr_comp g562 (.n_ena(w1084), .d(w29), .ena(w1085), .nres(w19), .nq(w226) );
	dmg_latchr_comp g563 (.n_ena(w191), .d(w16), .ena(w190), .nres(w19), .q(w1082), .nq(w1083) );
	dmg_latchr_comp g564 (.n_ena(w191), .d(w29), .ena(w190), .nres(w19), .q(w1106), .nq(w1105) );
	dmg_latchr_comp g565 (.n_ena(w191), .d(w55), .ena(w190), .nres(w19), .q(w1056), .nq(w847) );
	dmg_latchr_comp g566 (.n_ena(w191), .d(w187), .ena(w190), .nres(w19), .q(w1057), .nq(w1058) );
	dmg_latchr_comp g567 (.n_ena(w1089), .d(w16), .ena(w142), .nres(w1091), .nq(w310) );
	dmg_latchr_comp g568 (.n_ena(w1089), .d(w183), .ena(w142), .nres(w1091), .nq(w948) );
	dmg_latchr_comp g569 (.n_ena(w230), .d(w55), .ena(w142), .nres(w950), .nq(w949) );
	dmg_latchr_comp g570 (.n_ena(w952), .d(w55), .ena(w953), .nres(w954), .q(w23), .nq(w1112) );
	dmg_latchr_comp g571 (.n_ena(w669), .d(w55), .ena(w1134), .nres(w40), .q(w34), .nq(w35) );
	dmg_latchr_comp g572 (.n_ena(w669), .d(w187), .ena(w1134), .nres(w40), .q(w37), .nq(w36) );
	dmg_latchr_comp g573 (.n_ena(w380), .d(w589), .ena(w588), .nres(w523), .nq(w591) );
	dmg_latchr_comp g574 (.n_ena(w380), .d(w590), .ena(w381), .nres(w523), .nq(w524) );
	dmg_latchr_comp g575 (.n_ena(w520), .d(w578), .ena(w381), .nres(w523), .nq(w522) );
	dmg_latchr_comp g576 (.n_ena(w520), .d(w1174), .ena(w381), .nres(w523), .nq(w521) );
	dmg_nor g577 (.a(w90), .b(w3), .x(w2) );
	dmg_nor g578 (.a(w104), .b(w405), .x(w206) );
	dmg_not2 g579 (.a(w103), .x(w62) );
	dmg_nor g580 (.a(w110), .b(w1046), .x(w208) );
	dmg_nor g581 (.a(w761), .b(w416), .x(w967) );
	dmg_nor g582 (.a(w12), .b(w1108), .x(w13) );
	dmg_nor g583 (.a(w90), .b(w13), .x(w14) );
	dmg_nor g584 (.a(w550), .b(w70), .x(w1322) );
	dmg_nor g585 (.a(w70), .b(w1326), .x(w1329) );
	dmg_nor g586 (.a(w70), .b(w1054), .x(w1341) );
	dmg_nor g587 (.a(w70), .b(w1364), .x(w1325) );
	dmg_nor g588 (.a(w70), .b(w293), .x(w1146) );
	dmg_nor g589 (.a(w44), .b(w313), .x(w312) );
	dmg_nor g590 (.a(w1262), .b(w894), .x(w893) );
	dmg_nor g591 (.a(w1045), .b(w894), .x(w1044) );
	dmg_nor g592 (.a(w488), .b(w635), .x(w1315) );
	dmg_nor g593 (.a(w489), .b(w635), .x(w634) );
	dmg_nor g594 (.a(w489), .b(w636), .x(w490) );
	dmg_nor g595 (.a(w488), .b(w636), .x(w1314) );
	dmg_nor g596 (.a(w1050), .b(w894), .x(w831) );
	dmg_nor g597 (.a(w998), .b(w894), .x(w830) );
	dmg_nor g598 (.a(w456), .b(w61), .x(w60) );
	dmg_nor g599 (.a(w90), .b(w1135), .x(w89) );
	dmg_nor g600 (.a(w456), .b(w205), .x(w204) );
	dmg_nor g601 (.a(w90), .b(w1345), .x(w627) );
	dmg_not2 g602 (.a(w1259), .x(w399) );
	dmg_nor g603 (.a(w90), .b(w1251), .x(w1258) );
	dmg_nor g604 (.a(w1256), .b(w99), .x(w100) );
	dmg_nor g605 (.a(w348), .b(w664), .x(w108) );
	dmg_nor g606 (.a(w456), .b(w647), .x(w403) );
	dmg_nor g607 (.a(w456), .b(w404), .x(w210) );
	dmg_nor g608 (.a(w1338), .b(w70), .x(w1228) );
	dmg_nor g609 (.a(w768), .b(w416), .x(w1339) );
	dmg_nor g610 (.a(w767), .b(w416), .x(w417) );
	dmg_nor g611 (.a(w70), .b(w304), .x(w926) );
	dmg_nor g612 (.a(w168), .b(w27), .x(w161) );
	dmg_nor g613 (.a(w70), .b(w1128), .x(w1197) );
	dmg_nor g614 (.a(w70), .b(w876), .x(w877) );
	dmg_nor g615 (.a(w293), .b(w151), .x(w150) );
	dmg_nor g616 (.a(w70), .b(w144), .x(w145) );
	dmg_nor g617 (.a(w342), .b(w816), .x(w977) );
	dmg_nor g618 (.a(w146), .b(w162), .x(w147) );
	dmg_nor g619 (.a(w342), .b(w70), .x(w1077) );
	dmg_nor g620 (.a(w70), .b(w342), .x(w483) );
	dmg_nor g621 (.a(w342), .b(w272), .x(w136) );
	dmg_nor g622 (.a(w70), .b(w120), .x(w262) );
	dmg_nor g623 (.a(w984), .b(w70), .x(w1388) );
	dmg_nor g624 (.a(w532), .b(w70), .x(w476) );
	dmg_nor g625 (.a(w330), .b(w70), .x(w215) );
	dmg_nor g626 (.a(w726), .b(w456), .x(w457) );
	dmg_nor g627 (.a(w912), .b(w616), .x(w725) );
	dmg_nor g628 (.a(w913), .b(w175), .x(w176) );
	dmg_nor g629 (.a(w595), .b(w594), .x(w528) );
	dmg_nor g630 (.a(w596), .b(w597), .x(w655) );
	dmg_nor g631 (.a(w596), .b(w594), .x(w593) );
	dmg_nor g632 (.a(w70), .b(w251), .x(w270) );
	dmg_nor g633 (.a(w27), .b(w241), .x(w428) );
	dmg_nor g634 (.a(w241), .b(w240), .x(w239) );
	dmg_nor g635 (.a(w293), .b(w27), .x(w233) );
	dmg_nor g636 (.a(w70), .b(w238), .x(w216) );
	dmg_nor g637 (.a(w625), .b(w567), .x(w883) );
	dmg_nor g638 (.a(w369), .b(w370), .x(w1394) );
	dmg_nor g639 (.a(w564), .b(w567), .x(w565) );
	dmg_nor g640 (.a(w27), .b(w371), .x(w372) );
	dmg_nor g641 (.a(w1288), .b(w70), .x(w421) );
	dmg_nor g642 (.a(w1139), .b(w70), .x(w944) );
	dmg_nor g643 (.a(w853), .b(w567), .x(w568) );
	dmg_nor g644 (.a(w1395), .b(w567), .x(w946) );
	dmg_nor g645 (.a(w90), .b(w128), .x(w127) );
	dmg_nor g646 (.a(w1244), .b(w1138), .x(w1287) );
	dmg_nor g647 (.a(w1245), .b(w810), .x(w809) );
	dmg_nor g648 (.a(w692), .b(w691), .x(w609) );
	dmg_nor g649 (.a(w665), .b(w348), .x(w347) );
	dmg_nor g650 (.a(w349), .b(w70), .x(w95) );
	dmg_nor g651 (.a(w349), .b(w685), .x(w368) );
	dmg_nor g652 (.a(w369), .b(w686), .x(w678) );
	dmg_nor g653 (.a(w369), .b(w815), .x(w863) );
	dmg_nor g654 (.a(w70), .b(w1393), .x(w871) );
	dmg_nor g655 (.a(w70), .b(w798), .x(w792) );
	dmg_nor g656 (.a(w843), .b(w70), .x(w1375) );
	dmg_nor g657 (.a(w44), .b(w477), .x(w53) );
	dmg_nor g658 (.a(w70), .b(w71), .x(w860) );
	dmg_nor g659 (.a(w162), .b(w325), .x(w326) );
	dmg_nor g660 (.a(w533), .b(w70), .x(w324) );
	dmg_nor g661 (.a(w645), .b(w456), .x(w455) );
	dmg_nor g662 (.a(w410), .b(w70), .x(w346) );
	dmg_nor g663 (.a(w70), .b(w601), .x(w598) );
	dmg_nor g664 (.a(w70), .b(w605), .x(w604) );
	dmg_nor g665 (.a(w70), .b(w96), .x(w750) );
	dmg_nor g666 (.a(w70), .b(w748), .x(w1398) );
	dmg_nor g667 (.a(w456), .b(w1185), .x(w911) );
	dmg_nor g668 (.a(w456), .b(w1161), .x(w508) );
	dmg_nor g669 (.a(w507), .b(w456), .x(w505) );
	dmg_nor g670 (.a(w456), .b(w910), .x(w909) );
	dmg_nor g671 (.a(w1219), .b(w922), .x(w555) );
	dmg_nor g672 (.a(w35), .b(w37), .x(w1305) );
	dmg_nor g673 (.a(w34), .b(w37), .x(w33) );
	dmg_nor g674 (.a(w35), .b(w36), .x(w901) );
	dmg_nor g675 (.a(w34), .b(w36), .x(w895) );
	dmg_nor g676 (.a(w648), .b(w456), .x(w1311) );
	dmg_nor g677 (.a(w456), .b(w315), .x(w314) );
	dmg_nor g678 (.a(w456), .b(w64), .x(w65) );
	dmg_nor g679 (.a(w456), .b(w999), .x(w951) );
	dmg_nor g680 (.a(w970), .b(w894), .x(w1232) );
	dmg_nor g681 (.a(w66), .b(w67), .x(w345) );
	dmg_nor g682 (.a(w70), .b(w928), .x(w929) );
	dmg_nor g683 (.a(w293), .b(w27), .x(w292) );
	dmg_nor g684 (.a(w27), .b(w293), .x(w1036) );
	dmg_nor g685 (.a(w1035), .b(w147), .x(w148) );
	dmg_nor g686 (.a(w1145), .b(w70), .x(w308) );
	dmg_nor g687 (.a(w231), .b(w1098), .x(w1099) );
	dmg_nor g688 (.a(w70), .b(w1328), .x(w1007) );
	dmg_nor g689 (.a(w1360), .b(w70), .x(w1195) );
	dmg_nor g690 (.a(w1363), .b(w70), .x(w297) );
	dmg_nor g691 (.a(w44), .b(w1109), .x(w1108) );
	dmg_nor g692 (.a(w1213), .b(w1210), .x(w701) );
	dmg_nor g693 (.a(w1210), .b(w671), .x(w670) );
	dmg_nor g694 (.a(w90), .b(w700), .x(w628) );
	dmg_nor g695 (.a(w90), .b(w699), .x(w1049) );
	dmg_nor g696 (.a(w90), .b(w668), .x(w667) );
	dmg_nor g697 (.a(w395), .b(w396), .x(w397) );
	dmg_not3 g698 (.a(w1176), .x(w1175) );
	dmg_not3 g699 (.a(w1346), .x(w711) );
	dmg_not3 g700 (.a(w579), .x(w580) );
	dmg_not3 g701 (.a(w1096), .x(w1051) );
	dmg_not3 g702 (.a(w1090), .x(w231) );
	dmg_not3 g703 (.a(w1033), .x(w1200) );
	dmg_not3 g704 (.a(w1218), .x(w587) );
	dmg_not3 g705 (.a(w218), .x(w217) );
	dmg_not3 g706 (.a(w148), .x(w219) );
	dmg_not3 g707 (.a(w781), .x(w19) );
	dmg_not3 g708 (.a(w864), .x(w369) );
	dmg_not3 g709 (.a(w285), .x(w264) );
	dmg_not3 g710 (.a(w1321), .x(w1052) );
	dmg_not3 g711 (.a(w1318), .x(w1016) );
	dmg_not3 g712 (.a(w1309), .x(w965) );
	dmg_not2 g713 (.a(w14), .x(w15) );
	dmg_not2 g714 (.a(w142), .x(w1089) );
	dmg_not2 g715 (.a(w312), .x(w311) );
	dmg_not2 g716 (.a(w190), .x(w191) );
	dmg_not2 g717 (.a(w1108), .x(w225) );
	dmg_not2 g718 (.a(w996), .x(w1116) );
	dmg_not2 g719 (.a(w228), .x(w1115) );
	dmg_not2 g720 (.a(w656), .x(w657) );
	dmg_not2 g721 (.a(w1225), .x(w728) );
	dmg_not2 g722 (.a(w345), .x(w28) );
	dmg_not2 g723 (.a(w983), .x(w982) );
	dmg_not2 g724 (.a(w53), .x(w819) );
	dmg_not2 g725 (.a(w1193), .x(w243) );
	dmg_not2 g726 (.a(w440), .x(w780) );
	dmg_not2 g727 (.a(w1296), .x(w858) );
	dmg_not2 g728 (.a(w200), .x(w201) );
	dmg_not2 g729 (.a(w176), .x(w177) );
	dmg_not2 g730 (.a(w575), .x(w1142) );
	dmg_not2 g731 (.a(w1285), .x(w1391) );
	dmg_not2 g732 (.a(w817), .x(w339) );
	dmg_not2 g733 (.a(w725), .x(w530) );
	dmg_not2 g734 (.a(w208), .x(w646) );
	dmg_not2 g735 (.a(w317), .x(w316) );
	dmg_not2 g736 (.a(w62), .x(w63) );
	dmg_not2 g737 (.a(w209), .x(w207) );
	dmg_not2 g738 (.a(w673), .x(w209) );
	dmg_not2 g739 (.a(w296), .x(w162) );
	dmg_not2 g740 (.a(w70), .x(w1065) );
	dmg_not2 g741 (.a(w704), .x(w381) );
	dmg_not2 g742 (.a(w585), .x(w586) );
	dmg_not2 g743 (.a(w670), .x(w456) );
	dmg_not2 g744 (.a(w189), .x(w996) );
	dmg_not2 g745 (.a(w189), .x(w190) );
	dmg_not2 g746 (.a(w1095), .x(w285) );
	dmg_not2 g747 (.a(w1114), .x(w228) );
	dmg_not2 g748 (.a(w1114), .x(w1085) );
	dmg_not2 g749 (.a(w1085), .x(w1084) );
	dmg_nand g750 (.a(w188), .b(w204), .x(w1170) );
	dmg_nand g751 (.a(w180), .b(w295), .x(w1323) );
	dmg_nand g752 (.a(w1345), .b(w125), .x(w707) );
	dmg_nand g753 (.a(w1251), .b(w125), .x(w1257) );
	dmg_nand g754 (.a(w188), .b(w505), .x(w557) );
	dmg_nand g755 (.a(w1132), .b(w617), .x(w175) );
	dmg_nand g756 (.a(w55), .b(w30), .x(w562) );
	dmg_nand g757 (.a(w187), .b(w30), .x(w172) );
	dmg_nand g758 (.a(w637), .b(w508), .x(w514) );
	dmg_nand g759 (.a(w770), .b(w236), .x(w303) );
	dmg_nand g760 (.a(w881), .b(w236), .x(w265) );
	dmg_nand g761 (.a(w229), .b(w30), .x(w891) );
	dmg_nand g762 (.a(w183), .b(w30), .x(w1126) );
	dmg_nand g763 (.a(w180), .b(w30), .x(w795) );
	dmg_nand g764 (.a(w333), .b(w30), .x(w260) );
	dmg_nand g765 (.a(w505), .b(w504), .x(w503) );
	dmg_nand g766 (.a(w1349), .b(w643), .x(w1268) );
	dmg_nand g767 (.a(w338), .b(w42), .x(w916) );
	dmg_nand g768 (.a(w643), .b(w1406), .x(w47) );
	dmg_nand g769 (.a(w570), .b(w236), .x(w803) );
	dmg_nand g770 (.a(w255), .b(w236), .x(w254) );
	dmg_nand g771 (.a(w625), .b(w624), .x(w438) );
	dmg_nand g772 (.a(w564), .b(w624), .x(w884) );
	dmg_nand g773 (.a(w29), .b(w30), .x(w420) );
	dmg_nand g774 (.a(w16), .b(w30), .x(w1340) );
	dmg_nand g775 (.a(w853), .b(w624), .x(w945) );
	dmg_nand g776 (.a(w1395), .b(w624), .x(w947) );
	dmg_nand g777 (.a(w128), .b(w125), .x(w126) );
	dmg_nand g778 (.a(w1138), .b(w888), .x(w889) );
	dmg_nand g779 (.a(w810), .b(w624), .x(w811) );
	dmg_nand g780 (.a(w457), .b(w736), .x(w914) );
	dmg_nand g781 (.a(w643), .b(w188), .x(w1269) );
	dmg_nand g782 (.a(w508), .b(w1235), .x(w509) );
	dmg_nand g783 (.a(w571), .b(w234), .x(w1385) );
	dmg_nand g784 (.a(w796), .b(w234), .x(w235) );
	dmg_nand g785 (.a(w867), .b(w234), .x(w868) );
	dmg_nand g786 (.a(w827), .b(w617), .x(w616) );
	dmg_nand g787 (.a(w188), .b(w831), .x(w828) );
	dmg_nand g788 (.a(w637), .b(w505), .x(w541) );
	dmg_nand g789 (.a(w402), .b(w403), .x(w413) );
	dmg_nand g790 (.a(w643), .b(w402), .x(w401) );
	dmg_nand g791 (.a(w1135), .b(w125), .x(w1160) );
	dmg_nand g792 (.a(w188), .b(w1311), .x(w923) );
	dmg_nand g793 (.a(w188), .b(w65), .x(w1190) );
	dmg_nand g794 (.a(w1190), .b(w1138), .x(w30) );
	dmg_nand g795 (.a(w643), .b(w1188), .x(w1189) );
	dmg_nand g796 (.a(w188), .b(w951), .x(w1014) );
	dmg_nand g797 (.a(w1143), .b(w617), .x(w67) );
	dmg_nand g798 (.a(w637), .b(w831), .x(w69) );
	dmg_nand g799 (.a(w1005), .b(w941), .x(w1008) );
	dmg_nand g800 (.a(w643), .b(w836), .x(w835) );
	dmg_nand g801 (.a(w831), .b(w1103), .x(w1125) );
	dmg_nand g802 (.a(w831), .b(w1062), .x(w1061) );
	dmg_nand g803 (.a(w939), .b(w941), .x(w1087) );
	dmg_nand g804 (.a(w298), .b(w941), .x(w1199) );
	dmg_nand g805 (.a(w306), .b(w941), .x(w1320) );
	dmg_nand g806 (.a(w830), .b(w188), .x(w189) );
	dmg_nand g807 (.a(w333), .b(w295), .x(w305) );
	dmg_nand g808 (.a(w183), .b(w295), .x(w294) );
	dmg_nand g809 (.a(w951), .b(w1110), .x(w1113) );
	dmg_nand g810 (.a(w1044), .b(w188), .x(w1114) );
	dmg_nand g811 (.a(w637), .b(w951), .x(w952) );
	dmg_nand g812 (.a(w188), .b(w60), .x(w956) );
	dmg_nand g813 (.a(w414), .b(w60), .x(w415) );
	dmg_nand g814 (.a(w629), .b(w701), .x(w1218) );
	dmg_nand g815 (.a(w700), .b(w125), .x(w709) );
	dmg_nand g816 (.a(w699), .b(w125), .x(w1048) );
	dmg_nand g817 (.a(w188), .b(w643), .x(w715) );
	dmg_nand g818 (.a(w668), .b(w125), .x(w1263) );
	dmg_nand g819 (.a(w3), .b(w125), .x(w1157) );
	dmg_not6 g820 (.a(w389), .x(w390) );
	dmg_or g821 (.a(w90), .b(w1344), .x(w964) );
	dmg_or g822 (.a(w1099), .b(w231), .x(w1324) );
	dmg_or g823 (.a(w804), .b(w567), .x(w839) );
	dmg_or g824 (.a(w1078), .b(w1079), .x(w1075) );
	dmg_or g825 (.a(w70), .b(w342), .x(w987) );
	dmg_or g826 (.a(w620), .b(w621), .x(w1074) );
	dmg_or g827 (.a(w342), .b(w70), .x(w1193) );
	dmg_or g828 (.a(w1267), .b(w44), .x(w638) );
	dmg_or g829 (.a(w908), .b(w44), .x(w361) );
	dmg_or g830 (.a(w1220), .b(w93), .x(w94) );
	dmg_or g831 (.a(w1249), .b(w1142), .x(w781) );
	dmg_or g832 (.a(w778), .b(w472), .x(w427) );
	dmg_notif0 g833 (.n_ena(w225), .a(w1165), .x(w180) );
	dmg_notif0 g834 (.n_ena(w225), .a(w378), .x(w333) );
	dmg_notif0 g835 (.n_ena(w225), .a(w821), .x(w229) );
	dmg_notif0 g836 (.n_ena(w225), .a(w227), .x(w183) );
	dmg_notif0 g837 (.n_ena(w225), .a(w1163), .x(w16) );
	dmg_notif0 g838 (.n_ena(w225), .a(w1122), .x(w187) );
	dmg_notif0 g839 (.n_ena(w225), .a(w226), .x(w29) );
	dmg_notif0 g840 (.n_ena(w1061), .a(w995), .x(w183) );
	dmg_notif0 g841 (.n_ena(w311), .a(w948), .x(w183) );
	dmg_notif0 g842 (.n_ena(w311), .a(w1102), .x(w180) );
	dmg_notif0 g843 (.n_ena(w311), .a(w1092), .x(w333) );
	dmg_notif0 g844 (.n_ena(w311), .a(w949), .x(w55) );
	dmg_notif0 g845 (.n_ena(w311), .a(w1090), .x(w229) );
	dmg_notif0 g846 (.n_ena(w311), .a(w1086), .x(w29) );
	dmg_notif0 g847 (.n_ena(w311), .a(w310), .x(w16) );
	dmg_notif0 g848 (.n_ena(w15), .a(w20), .x(w183) );
	dmg_notif0 g849 (.n_ena(w15), .a(w20), .x(w16) );
	dmg_notif0 g850 (.n_ena(w15), .a(w20), .x(w180) );
	dmg_notif0 g851 (.n_ena(w15), .a(w20), .x(w229) );
	dmg_notif0 g852 (.n_ena(w15), .a(w20), .x(w333) );
	dmg_notif0 g853 (.n_ena(w15), .a(w20), .x(w55) );
	dmg_notif0 g854 (.n_ena(w649), .a(w35), .x(w55) );
	dmg_notif0 g855 (.n_ena(w649), .a(w36), .x(w187) );
	dmg_notif0 g856 (.n_ena(w415), .a(w636), .x(w187) );
	dmg_notif0 g857 (.n_ena(w1001), .a(w1002), .x(w180) );
	dmg_notif0 g858 (.n_ena(w1001), .a(w1131), .x(w333) );
	dmg_notif0 g859 (.n_ena(w116), .a(w804), .x(w16) );
	dmg_notif0 g860 (.n_ena(w819), .a(w1105), .x(w29) );
	dmg_notif0 g861 (.n_ena(w819), .a(w847), .x(w55) );
	dmg_notif0 g862 (.n_ena(w835), .a(w834), .x(w183) );
	dmg_notif0 g863 (.n_ena(w819), .a(w1058), .x(w187) );
	dmg_notif0 g864 (.n_ena(w819), .a(w1083), .x(w16) );
	dmg_notif0 g865 (.n_ena(w1125), .a(w77), .x(w55) );
	dmg_notif0 g866 (.n_ena(w819), .a(w824), .x(w180) );
	dmg_notif0 g867 (.n_ena(w819), .a(w1117), .x(w333) );
	dmg_notif0 g868 (.n_ena(w1189), .a(w973), .x(w333) );
	dmg_notif0 g869 (.n_ena(w552), .a(w745), .x(w55) );
	dmg_notif0 g870 (.n_ena(w530), .a(w1335), .x(w16) );
	dmg_notif0 g871 (.n_ena(w530), .a(w1337), .x(w29) );
	dmg_notif0 g872 (.n_ena(w530), .a(w529), .x(w187) );
	dmg_notif0 g873 (.n_ena(w361), .a(w360), .x(w229) );
	dmg_notif0 g874 (.n_ena(w413), .a(w412), .x(w187) );
	dmg_notif0 g875 (.n_ena(w509), .a(w510), .x(w55) );
	dmg_notif0 g876 (.n_ena(w28), .a(w1203), .x(w55) );
	dmg_notif0 g877 (.n_ena(w28), .a(w539), .x(w16) );
	dmg_notif0 g878 (.n_ena(w28), .a(w331), .x(w333) );
	dmg_notif0 g879 (.n_ena(w478), .a(w979), .x(w29) );
	dmg_notif0 g880 (.n_ena(w478), .a(w1123), .x(w55) );
	dmg_notif0 g881 (.n_ena(w478), .a(w980), .x(w16) );
	dmg_notif0 g882 (.n_ena(w487), .a(w1384), .x(w16) );
	dmg_notif0 g883 (.n_ena(w487), .a(w622), .x(w229) );
	dmg_notif0 g884 (.n_ena(w116), .a(w786), .x(w229) );
	dmg_notif0 g885 (.n_ena(w435), .a(w434), .x(w187) );
	dmg_notif0 g886 (.n_ena(w212), .a(w1297), .x(w333) );
	dmg_notif0 g887 (.n_ena(w212), .a(w1242), .x(w183) );
	dmg_notif0 g888 (.n_ena(w212), .a(w376), .x(w180) );
	dmg_notif0 g889 (.n_ena(w177), .a(w465), .x(w229) );
	dmg_notif0 g890 (.n_ena(w177), .a(w640), .x(w183) );
	dmg_notif0 g891 (.n_ena(w177), .a(w642), .x(w16) );
	dmg_notif0 g892 (.n_ena(w615), .a(w1365), .x(w333) );
	dmg_notif0 g893 (.n_ena(w615), .a(w614), .x(w180) );
	dmg_notif0 g894 (.n_ena(w177), .a(w192), .x(w29) );
	dmg_notif0 g895 (.n_ena(w174), .a(w1301), .x(w333) );
	dmg_notif0 g896 (.n_ena(w174), .a(w184), .x(w183) );
	dmg_notif0 g897 (.n_ena(w177), .a(w186), .x(w187) );
	dmg_notif0 g898 (.n_ena(w177), .a(w462), .x(w55) );
	dmg_notif0 g899 (.n_ena(w177), .a(w450), .x(w333) );
	dmg_notif0 g900 (.n_ena(w177), .a(w178), .x(w180) );
	dmg_notif0 g901 (.n_ena(w116), .a(w626), .x(w29) );
	dmg_notif0 g902 (.n_ena(w28), .a(w1140), .x(w29) );
	dmg_notif0 g903 (.n_ena(w28), .a(w257), .x(w229) );
	dmg_notif0 g904 (.n_ena(w28), .a(w573), .x(w180) );
	dmg_notif0 g905 (.n_ena(w116), .a(w783), .x(w183) );
	dmg_notif0 g906 (.n_ena(w116), .a(w117), .x(w180) );
	dmg_notif0 g907 (.n_ena(w916), .a(w789), .x(w229) );
	dmg_notif0 g908 (.n_ena(w46), .a(w138), .x(w183) );
	dmg_notif0 g909 (.n_ena(w46), .a(w334), .x(w333) );
	dmg_notif0 g910 (.n_ena(w46), .a(w1286), .x(w180) );
	dmg_notif0 g911 (.n_ena(w47), .a(w1020), .x(w229) );
	dmg_notif0 g912 (.n_ena(w487), .a(w54), .x(w55) );
	dmg_notif0 g913 (.n_ena(w487), .a(w486), .x(w187) );
	dmg_notif0 g914 (.n_ena(w487), .a(w1284), .x(w29) );
	dmg_notif0 g915 (.n_ena(w478), .a(w479), .x(w187) );
	dmg_notif0 g916 (.n_ena(w435), .a(w436), .x(w229) );
	dmg_notif0 g917 (.n_ena(w435), .a(w856), .x(w55) );
	dmg_notif0 g918 (.n_ena(w435), .a(w857), .x(w29) );
	dmg_notif0 g919 (.n_ena(w503), .a(w502), .x(w55) );
	dmg_notif0 g920 (.n_ena(w435), .a(w213), .x(w16) );
	dmg_notif0 g921 (.n_ena(w1268), .a(w1249), .x(w187) );
	dmg_notif0 g922 (.n_ena(w361), .a(w352), .x(w16) );
	dmg_notif0 g923 (.n_ena(w361), .a(w351), .x(w55) );
	dmg_notif0 g924 (.n_ena(w361), .a(w561), .x(w29) );
	dmg_notif0 g925 (.n_ena(w361), .a(w362), .x(w187) );
	dmg_notif0 g926 (.n_ena(w638), .a(w735), .x(w183) );
	dmg_notif0 g927 (.n_ena(w638), .a(w366), .x(w333) );
	dmg_notif0 g928 (.n_ena(w638), .a(w639), .x(w180) );
	dmg_notif0 g929 (.n_ena(w914), .a(w594), .x(w16) );
	dmg_notif0 g930 (.n_ena(w914), .a(w596), .x(w55) );
	dmg_notif0 g931 (.n_ena(w615), .a(w915), .x(w183) );
	dmg_notif0 g932 (.n_ena(w174), .a(w1272), .x(w180) );
	dmg_notif0 g933 (.n_ena(w559), .a(w1276), .x(w183) );
	dmg_notif0 g934 (.n_ena(w559), .a(w660), .x(w29) );
	dmg_notif0 g935 (.n_ena(w559), .a(w675), .x(w333) );
	dmg_notif0 g936 (.n_ena(w559), .a(w107), .x(w180) );
	dmg_notif0 g937 (.n_ena(w552), .a(w753), .x(w183) );
	dmg_notif0 g938 (.n_ena(w559), .a(w106), .x(w229) );
	dmg_notif0 g939 (.n_ena(w552), .a(w1226), .x(w229) );
	dmg_notif0 g940 (.n_ena(w552), .a(w746), .x(w333) );
	dmg_notif0 g941 (.n_ena(w552), .a(w1254), .x(w180) );
	dmg_notif0 g942 (.n_ena(w401), .a(w400), .x(w180) );
	dmg_notif0 g943 (.n_ena(w28), .a(w919), .x(w187) );
	dmg_notif0 g944 (.n_ena(w28), .a(w328), .x(w183) );
	dmg_notif0 g945 (.n_ena(w68), .a(w1013), .x(w333) );
	dmg_notif0 g946 (.n_ena(w68), .a(w832), .x(w180) );
	dmg_notif0 g947 (.n_ena(w68), .a(w918), .x(w183) );
	dmg_notif0 g948 (.n_ena(w1001), .a(w975), .x(w183) );
	dmg_notif0 g949 (.n_ena(w415), .a(w488), .x(w55) );
	dmg_notif0 g950 (.n_ena(w1113), .a(w1112), .x(w55) );
	dmg_notif0 g951 (.n_ena(w15), .a(w20), .x(w29) );
	dmg_notif0 g952 (.n_ena(w15), .a(w20), .x(w187) );
	dmg_notif0 g953 (.n_ena(w819), .a(w1166), .x(w183) );
	dmg_notif0 g954 (.n_ena(w819), .a(w820), .x(w229) );
	dmg_notif0 g955 (.n_ena(w225), .a(w224), .x(w55) );
	dmg_and g956 (.a(w1071), .b(w132), .x(w131) );
	dmg_and g957 (.a(w133), .b(w132), .x(w1081) );
	dmg_and g958 (.a(w941), .b(w1327), .x(w1326) );
	dmg_and g959 (.a(w941), .b(w1053), .x(w1054) );
	dmg_and g960 (.a(w156), .b(w155), .x(w549) );
	dmg_and g961 (.a(w443), .b(w475), .x(w548) );
	dmg_and g962 (.a(w545), .b(w475), .x(w547) );
	dmg_and g963 (.a(w474), .b(w475), .x(w546) );
	dmg_and g964 (.a(w295), .b(w551), .x(w550) );
	dmg_and g965 (.a(w295), .b(w1361), .x(w1360) );
	dmg_and g966 (.a(w357), .b(w356), .x(w1359) );
	dmg_and g967 (.a(w1222), .b(w356), .x(w1358) );
	dmg_and g968 (.a(w355), .b(w356), .x(w1357) );
	dmg_and g969 (.a(w91), .b(w356), .x(w1342) );
	dmg_and g970 (.a(w1214), .b(w188), .x(w637) );
	dmg_and g971 (.a(w1356), .b(w887), .x(w808) );
	dmg_and g972 (.a(w719), .b(w805), .x(w1047) );
	dmg_and g973 (.a(w188), .b(w60), .x(w630) );
	dmg_and g974 (.a(w932), .b(w933), .x(w1280) );
	dmg_and g975 (.a(w24), .b(w23), .x(w22) );
	dmg_and g976 (.a(w833), .b(w921), .x(w154) );
	dmg_and g977 (.a(w188), .b(w314), .x(w142) );
	dmg_and g978 (.a(w838), .b(w837), .x(w1062) );
	dmg_and g979 (.a(w845), .b(w272), .x(w994) );
	dmg_and g980 (.a(w223), .b(w617), .x(w618) );
	dmg_and g981 (.a(w76), .b(w75), .x(w1080) );
	dmg_and g982 (.a(w236), .b(w880), .x(w876) );
	dmg_and g983 (.a(w236), .b(w974), .x(w1128) );
	dmg_and g984 (.a(w30), .b(w769), .x(w768) );
	dmg_and g985 (.a(w30), .b(w516), .x(w767) );
	dmg_and g986 (.a(w491), .b(w492), .x(w497) );
	dmg_and g987 (.a(w497), .b(w496), .x(w633) );
	dmg_and g988 (.a(w30), .b(w31), .x(w1338) );
	dmg_and g989 (.a(w319), .b(w318), .x(w42) );
	dmg_and g990 (.a(w32), .b(w902), .x(w903) );
	dmg_and g991 (.a(w909), .b(w188), .x(w1225) );
	dmg_and g992 (.a(w911), .b(w188), .x(w1265) );
	dmg_and g993 (.a(w29), .b(w90), .x(w1266) );
	dmg_and g994 (.a(w188), .b(w643), .x(w644) );
	dmg_and g995 (.a(w188), .b(w909), .x(w680) );
	dmg_and g996 (.a(w500), .b(w501), .x(w1207) );
	dmg_and g997 (.a(w403), .b(w188), .x(w1206) );
	dmg_and g998 (.a(w210), .b(w188), .x(w1296) );
	dmg_and g999 (.a(w893), .b(w188), .x(w817) );
	dmg_and g1000 (.a(w188), .b(w42), .x(w983) );
	dmg_and g1001 (.a(w1019), .b(w482), .x(w1018) );
	dmg_and g1002 (.a(w234), .b(w797), .x(w798) );
	dmg_and g1003 (.a(w234), .b(w799), .x(w1393) );
	dmg_and g1004 (.a(w455), .b(w188), .x(w200) );
	dmg_and g1005 (.a(w508), .b(w188), .x(w454) );
	dmg_and g1006 (.a(w455), .b(w188), .x(w203) );
	dmg_and g1007 (.a(w30), .b(w469), .x(w1288) );
	dmg_and g1008 (.a(w30), .b(w1246), .x(w1139) );
	dmg_and g1009 (.a(w234), .b(w271), .x(w251) );
	dmg_and g1010 (.a(w236), .b(w872), .x(w238) );
	dmg_and g1011 (.a(w236), .b(w237), .x(w240) );
	dmg_and g1012 (.a(w188), .b(w42), .x(w1285) );
	dmg_and g1013 (.a(w188), .b(w210), .x(w730) );
	dmg_and g1014 (.a(w188), .b(w457), .x(w1369) );
	dmg_and g1015 (.a(w505), .b(w188), .x(w181) );
	dmg_and g1016 (.a(w1273), .b(w692), .x(w603) );
	dmg_and g1017 (.a(w664), .b(w665), .x(w661) );
	dmg_and g1018 (.a(w1255), .b(w1256), .x(w676) );
	dmg_and g1019 (.a(w30), .b(w531), .x(w532) );
	dmg_and g1020 (.a(w30), .b(w1196), .x(w984) );
	dmg_and g1021 (.a(w30), .b(w329), .x(w330) );
	dmg_and g1022 (.a(w76), .b(w617), .x(w838) );
	dmg_and g1023 (.a(w166), .b(w162), .x(w163) );
	dmg_and g1024 (.a(w188), .b(w951), .x(w295) );
	dmg_and g1025 (.a(w188), .b(w893), .x(w1191) );
	dmg_and g1026 (.a(w766), .b(w512), .x(w511) );
	dmg_and g1027 (.a(w896), .b(w899), .x(w32) );
	dmg_and g1028 (.a(w319), .b(w320), .x(w643) );
	dmg_and g1029 (.a(w592), .b(w528), .x(w721) );
	dmg_and g1030 (.a(w399), .b(w653), .x(w760) );
	dmg_and g1031 (.a(w399), .b(w722), .x(w1348) );
	dmg_and g1032 (.a(w399), .b(w723), .x(w1046) );
	dmg_and g1033 (.a(w399), .b(w721), .x(w720) );
	dmg_and g1034 (.a(w188), .b(w204), .x(w1134) );
	dmg_and g1035 (.a(w188), .b(w701), .x(w579) );
	dmg_and g1036 (.a(w295), .b(w1362), .x(w1363) );
	dmg_and g1037 (.a(w941), .b(w1006), .x(w1328) );
	dmg_and g1038 (.a(w1100), .b(w1101), .x(w259) );
	dmg_and g1039 (.a(w129), .b(w132), .x(w130) );
	dmg_and g1040 (.a(w841), .b(w132), .x(w1164) );
	dmg_nand4 g1041 (.a(w1216), .b(w1212), .c(w583), .d(w111), .x(w1213) );
	dmg_nand4 g1042 (.a(w959), .b(w113), .c(w807), .d(w808), .x(w574) );
	dmg_nand4 g1043 (.a(w207), .b(w62), .c(w316), .d(w646), .x(w645) );
	dmg_nand4 g1044 (.a(w208), .b(w316), .c(w62), .d(w209), .x(w999) );
	dmg_nand4 g1045 (.a(w209), .b(w63), .c(w316), .d(w646), .x(w507) );
	dmg_nand4 g1046 (.a(w646), .b(w206), .c(w63), .d(w209), .x(w647) );
	dmg_nand4 g1047 (.a(w207), .b(w63), .c(w206), .d(w646), .x(w648) );
	dmg_nand4 g1048 (.a(w208), .b(w206), .c(w63), .d(w207), .x(w64) );
	dmg_nand4 g1049 (.a(w209), .b(w62), .c(w316), .d(w646), .x(w726) );
	dmg_nand4 g1050 (.a(w209), .b(w62), .c(w316), .d(w208), .x(w1045) );
	dmg_nand4 g1051 (.a(w208), .b(w206), .c(w62), .d(w209), .x(w315) );
	dmg_nand4 g1052 (.a(w208), .b(w206), .c(w63), .d(w209), .x(w404) );
	dmg_nand4 g1053 (.a(w208), .b(w316), .c(w63), .d(w209), .x(w205) );
	dmg_nand4 g1054 (.a(w207), .b(w63), .c(w206), .d(w208), .x(w1050) );
	dmg_nand4 g1055 (.a(w646), .b(w206), .c(w62), .d(w207), .x(w1161) );
	dmg_nand4 g1056 (.a(w207), .b(w62), .c(w206), .d(w208), .x(w1262) );
	dmg_nand4 g1057 (.a(w208), .b(w206), .c(w62), .d(w207), .x(w61) );
	dmg_nand4 g1058 (.a(w207), .b(w62), .c(w316), .d(w208), .x(w998) );
	dmg_nand4 g1059 (.a(w208), .b(w316), .c(w63), .d(w207), .x(w910) );
	dmg_nand4 g1060 (.a(w646), .b(w206), .c(w62), .d(w209), .x(w1185) );
	dmg_nand4 g1061 (.a(w209), .b(w62), .c(w206), .d(w208), .x(w970) );
	dmg_mux g1062 (.sel(w399), .d1(w102), .d0(w103), .q(w1354) );
	dmg_mux g1063 (.sel(w399), .d1(w105), .d0(w104), .q(w1154) );
	dmg_mux g1064 (.sel(w399), .d1(w109), .d0(w110), .q(w1155) );
	dmg_mux g1065 (.sel(w399), .d1(w398), .d0(w713), .q(w1176) );
	dmg_mux g1066 (.sel(w385), .d1(w383), .d0(w384), .q(w1345) );
	dmg_mux g1067 (.sel(w385), .d1(w581), .d0(w582), .q(w1251) );
	dmg_mux g1068 (.sel(w385), .d1(w1355), .d0(w4), .q(w3) );
	dmg_mux g1069 (.sel(w385), .d1(w1137), .d0(w1136), .q(w668) );
	dmg_mux g1070 (.sel(w385), .d1(w387), .d0(w386), .q(w1135) );
	dmg_mux g1071 (.sel(w385), .d1(w697), .d0(w698), .q(w699) );
	dmg_mux g1072 (.sel(w385), .d1(w584), .d0(w696), .q(w700) );
	dmg_mux g1073 (.sel(w385), .d1(w7), .d0(w6), .q(w128) );
	dmg_mux g1074 (.sel(w838), .d1(w480), .d0(w1018), .q(w619) );
	dmg_mux g1075 (.sel(w1038), .d1(w141), .d0(w264), .q(w865) );
	dmg_mux g1076 (.sel(w981), .d1(w1076), .d0(w1075), .q(w480) );
	dmg_mux g1077 (.sel(w1038), .d1(w141), .d0(w1200), .q(w1319) );
	dmg_mux g1078 (.sel(w1038), .d1(w141), .d0(w1051), .q(w1310) );
	dmg_mux g1079 (.sel(w399), .d1(w588), .d0(w587), .q(w1346) );
	dmg_mux g1080 (.sel(w399), .d1(w674), .d0(w673), .q(w1153) );
	dmg_bufif0 g1081 (.a0(w1158), .n_ena(w125), .a1(w1158), .x(w104) );
	dmg_bufif0 g1082 (.a0(w124), .n_ena(w125), .a1(w124), .x(w111) );
	dmg_bufif0 g1083 (.a0(w695), .n_ena(w125), .a1(w695), .x(w110) );
	dmg_bufif0 g1084 (.a0(w1173), .n_ena(w125), .a1(w1173), .x(w583) );
	dmg_bufif0 g1085 (.a0(w87), .n_ena(w125), .a1(w87), .x(w672) );
	dmg_bufif0 g1086 (.a0(w997), .n_ena(w125), .a1(w997), .x(w112) );
	dmg_bufif0 g1087 (.a0(w705), .n_ena(w125), .a1(w705), .x(w103) );
	dmg_nor_latch g1088 (.s(w739), .r(w689), .q(w688) );
	dmg_nor_latch g1089 (.s(w569), .r(w429), .q(w430) );
	dmg_nor_latch g1090 (.s(w861), .r(w120), .nq(w862) );
	dmg_nor_latch g1091 (.s(w342), .r(w844), .q(w1019) );
	dmg_nor_latch g1092 (.s(w1281), .r(w987), .q(w986) );
	dmg_nor_latch g1093 (.s(w925), .r(w928), .nq(w927) );
	dmg_nor_latch g1094 (.s(w348), .r(w409), .q(w408) );
	dmg_nor_latch g1095 (.s(w744), .r(w601), .nq(w743) );
	dmg_nor_latch g1096 (.s(w751), .r(w748), .nq(w749) );
	dmg_nor_latch g1097 (.s(w922), .r(w931), .q(w932) );
	dmg_nor_latch g1098 (.s(w27), .r(w1317), .q(w833) );
	dmg_bufif0 g1099 (.a0(w446), .n_ena(w125), .a1(w446), .x(w673) );
	dmg_not2 g1100 (.a(w397), .x(w398) );
	dmg_latch g1101 (.ena(w5), .d(w103), .q(w384) );
	dmg_latch g1102 (.ena(w5), .d(w583), .q(w4) );
	dmg_latch g1103 (.ena(w5), .d(w112), .q(w582) );
	dmg_latch g1104 (.ena(w5), .d(w110), .q(w1136) );
	dmg_latch g1105 (.ena(w5), .d(w672), .q(w386) );
	dmg_latch g1106 (.ena(w5), .d(w111), .q(w696) );
	dmg_latch g1107 (.ena(w5), .d(w673), .q(w6) );
	dmg_latch g1108 (.ena(w5), .d(w104), .q(w698) );
	dmg_latch g1109 (.ena(w10), .d(w886), .q(w1215) );
	dmg_latch g1110 (.ena(w116), .d(w788), .q(w117) );
	dmg_latch g1111 (.ena(w116), .d(w784), .q(w783) );
	dmg_latch g1112 (.ena(w116), .d(w785), .q(w439) );
	dmg_latch g1113 (.ena(w116), .d(w787), .q(w786) );
	dmg_not4 g1114 (.a(w143), .x(w144) );
	dmg_dffsr g1115 (.nset1(w1087), .nset2(w1087), .d(w307), .q(w1088), .nres(w1325), .clk(w1052) );
	dmg_dffsr g1116 (.nset1(w305), .nset2(w305), .d(w1041), .q(w939), .nres(w1195), .clk(w1042) );
	dmg_dffsr g1117 (.nset1(w891), .nset2(w891), .d(w890), .q(w570), .nres(w1388), .clk(w259) );
	dmg_dffsr g1118 (.nset1(w1008), .nset2(w1008), .d(w1009), .q(w302), .nres(w1007), .clk(w1052) );
	dmg_dffsr g1119 (.nset1(w1199), .nset2(w1199), .d(w1088), .q(w1009), .nres(w1341), .clk(w1052) );
	dmg_dffsr g1120 (.nset1(w1385), .nset2(w1385), .d(w801), .q(w800), .nres(w871), .clk(w219) );
	dmg_dffsr g1121 (.nset1(w260), .nset2(w260), .d(w812), .q(w796), .nres(w215), .clk(w259) );
	dmg_dffsr g1122 (.nset1(w254), .nset2(w254), .d(w878), .q(w232), .nres(w216), .clk(w217) );
	dmg_dffsr g1123 (.nset1(w803), .nset2(w803), .d(w232), .q(w801), .nres(w239), .clk(w217) );
	dmg_dffsr g1124 (.nset1(w235), .nset2(w235), .d(w800), .q(w869), .nres(w792), .clk(w219) );
	dmg_dffsr g1125 (.nset1(w562), .nset2(w562), .d(w1230), .q(w770), .nres(w1228), .clk(w259) );
	dmg_dffsr g1126 (.nset1(w172), .nset2(w172), .d(w1141), .q(w1005), .nres(w1339), .clk(w259) );
	dmg_dffsr g1127 (.nset1(w795), .nset2(w795), .d(w794), .q(w571), .nres(w476), .clk(w259) );
	dmg_dffsr g1128 (.nset1(w1340), .nset2(w1340), .d(w775), .q(w881), .nres(w944), .clk(w259) );
	dmg_dffsr g1129 (.nset1(w1126), .nset2(w1126), .d(w418), .q(w867), .nres(w417), .clk(w259) );
	dmg_dffsr g1130 (.nset1(w868), .nset2(w868), .d(w869), .q(w269), .nres(w270), .clk(w219) );
	dmg_dffsr g1131 (.nset1(w265), .nset2(w265), .d(w266), .q(w878), .nres(w877), .clk(w217) );
	dmg_dffsr g1132 (.nset1(w303), .nset2(w303), .d(w302), .q(w266), .nres(w1197), .clk(w217) );
	dmg_dffsr g1133 (.nset1(w420), .nset2(w420), .d(w422), .q(w255), .nres(w421), .clk(w259) );
	dmg_dffsr g1134 (.nset1(w294), .nset2(w294), .d(w1012), .q(w298), .nres(w297), .clk(w1042) );
	dmg_dffsr g1135 (.nset1(w1320), .nset2(w1320), .d(w20), .q(w307), .nres(w1329), .clk(w1052) );
	dmg_not6 g1136 (.a(w44), .x(w629) );
	dmg_not6 g1137 (.a(w712), .x(w713) );
	dmg_mux g1138 (.sel(w617), .d1(w85), .d0(w965), .q(w84) );
	dmg_not6 g1139 (.a(w806), .x(w188) );
	dmg_not6 g1140 (.a(w1223), .x(w1224) );
	dmg_not6 g1141 (.a(w782), .x(w241) );
	dmg_dffr_comp g1142 (.nr1(w780), .nr2(w780), .d(w267), .ck(w144), .cck(w779), .q(w253) );
	dmg_dffr_comp g1143 (.nr1(w299), .nr2(w299), .d(w796), .ck(w144), .cck(w471), .q(w426) );
	dmg_dffr_comp g1144 (.nr1(w299), .nr2(w299), .d(w882), .ck(w144), .cck(w774), .q(w1403) );
	dmg_dffr_comp g1145 (.nr1(w299), .nr2(w299), .d(w570), .ck(w144), .cck(w471), .q(w252) );
	dmg_dffr_comp g1146 (.nr1(w299), .nr2(w299), .d(w255), .ck(w144), .cck(w771), .q(w777) );
	dmg_dffr_comp g1147 (.nr1(w299), .nr2(w299), .d(w867), .ck(w144), .cck(w471), .q(w942) );
	dmg_dffr_comp g1148 (.nr1(w299), .nr2(w299), .d(w419), .ck(w144), .cck(w774), .q(w773) );
	dmg_dffr_comp g1149 (.nr1(w299), .nr2(w299), .d(w875), .ck(w144), .cck(w300), .q(w873) );
	dmg_dffr_comp g1150 (.nr1(w299), .nr2(w299), .d(w943), .ck(w144), .cck(w300), .q(w879) );
	dmg_dffr_comp g1151 (.nr1(w299), .nr2(w299), .d(w301), .ck(w144), .cck(w300), .q(w936) );
	dmg_dffr_comp g1152 (.nr1(w299), .nr2(w299), .d(w770), .ck(w144), .cck(w938), .q(w1039) );
	dmg_dffr_comp g1153 (.nr1(w299), .nr2(w299), .d(w1144), .ck(w144), .cck(w300), .q(w935) );
	dmg_dffr_comp g1154 (.nr1(w299), .nr2(w299), .d(w939), .ck(w144), .cck(w938), .q(w874) );
	dmg_dffr_comp g1155 (.nr1(w780), .nr2(w780), .d(w268), .ck(w144), .cck(w779), .q(w814) );
	dmg_dffr_comp g1156 (.nr1(w780), .nr2(w780), .d(w870), .ck(w144), .cck(w779), .q(w793) );
	dmg_dffr_comp g1157 (.nr1(w780), .nr2(w780), .d(w866), .ck(w144), .cck(w779), .q(w802) );
	dmg_dffr_comp g1158 (.nr1(w299), .nr2(w299), .d(w571), .ck(w144), .cck(w471), .q(w470) );
	dmg_dffr_comp g1159 (.nr1(w299), .nr2(w299), .d(w306), .ck(w144), .cck(w771), .q(w1400) );
	dmg_dffr_comp g1160 (.nr1(w299), .nr2(w299), .d(w1005), .ck(w144), .cck(w938), .q(w937) );
	dmg_dffr_comp g1161 (.nr1(w299), .nr2(w299), .d(w1010), .ck(w144), .cck(w774), .q(w1399) );
	dmg_dffr_comp g1162 (.nr1(w299), .nr2(w299), .d(w298), .ck(w144), .cck(w938), .q(w934) );
	dmg_not4 g1163 (.a(w123), .x(w122) );
	dmg_dffr_comp g1164 (.nr1(w299), .nr2(w299), .d(w881), .ck(w144), .cck(w771), .q(w772) );
	dmg_or g1165 (.a(w45), .b(w44), .x(w46) );
	dmg_or g1166 (.a(w43), .b(w44), .x(w478) );
	dmg_or g1167 (.a(w1376), .b(w1377), .x(w48) );
	dmg_or g1168 (.a(w241), .b(w27), .x(w440) );
	dmg_or g1169 (.a(w241), .b(w27), .x(w429) );
	dmg_or g1170 (.a(w626), .b(w567), .x(w566) );
	dmg_or g1171 (.a(w1234), .b(w44), .x(w435) );
	dmg_or g1172 (.a(w211), .b(w44), .x(w212) );
	dmg_or g1173 (.a(w727), .b(w616), .x(w615) );
	dmg_or g1174 (.a(w70), .b(w349), .x(w689) );
	dmg_or g1175 (.a(w1353), .b(w175), .x(w174) );
	dmg_or g1176 (.a(w1000), .b(w67), .x(w68) );
	dmg_or g1177 (.a(w619), .b(w618), .x(w132) );
	dmg_or g1178 (.a(w154), .b(w617), .x(w155) );
	dmg_or g1179 (.a(w1280), .b(w617), .x(w356) );
	dmg_or g1180 (.a(w1111), .b(w44), .x(w1001) );
	dmg_or g1181 (.a(w1209), .b(w1210), .x(w894) );
	dmg_aon22 g1182 (.a0(w134), .a1(w1071), .b0(w1282), .b1(w622), .x(w1072) );
	dmg_aon22 g1183 (.a0(w134), .a1(w129), .b0(w1070), .b1(w622), .x(w1073) );
	dmg_aon22 g1184 (.a0(w134), .a1(w133), .b0(w988), .b1(w622), .x(w842) );
	dmg_aon22 g1185 (.a0(w1221), .a1(w679), .b0(w679), .b1(w360), .x(w907) );
	dmg_aon22 g1186 (.a0(w1221), .a1(w355), .b0(w906), .b1(w360), .x(w905) );
	dmg_aon22 g1187 (.a0(w506), .a1(w91), .b0(w904), .b1(w360), .x(w359) );
	dmg_aon22 g1188 (.a0(w506), .a1(w357), .b0(w358), .b1(w360), .x(w364) );
	dmg_aon22 g1189 (.a0(w654), .a1(w528), .b0(w592), .b1(w655), .x(w723) );
	dmg_aon22 g1190 (.a0(w442), .a1(w443), .b0(w444), .b1(w436), .x(w535) );
	dmg_aon22 g1191 (.a0(w442), .a1(w437), .b0(w437), .b1(w436), .x(w445) );
	dmg_aon22 g1192 (.a0(w442), .a1(w545), .b0(w537), .b1(w436), .x(w854) );
	dmg_aon22 g1193 (.a0(w442), .a1(w156), .b0(w536), .b1(w436), .x(w157) );
	dmg_aon22 g1194 (.a0(w51), .a1(w790), .b0(w789), .b1(w791), .x(w247) );
	dmg_muxi g1195 (.sel(w525), .d1(w522), .d0(w521), .q(w654) );
	dmg_muxi g1196 (.sel(w525), .d1(w524), .d0(w591), .q(w592) );
	dmg_muxi g1197 (.sel(w624), .d1(w56), .d0(w57), .q(w1247) );
	dmg_muxi g1198 (.sel(w525), .d1(w526), .d0(w1261), .q(w527) );
	dmg_muxi g1199 (.sel(w525), .d1(w757), .d0(w758), .q(w724) );
	dmg_nand_latch g1200 (.nr(w346), .ns(w690), .nq(w691) );
	dmg_nand_latch g1201 (.nr(w145), .ns(w150), .nq(w146) );
	dmg_nand_latch g1202 (.nr(w1375), .ns(w1374), .nq(w1376) );
	dmg_nand_latch g1203 (.nr(w967), .ns(w98), .nq(w99) );
	dmg_not g1204 (.a(w557), .x(w558) );
	dmg_nand g1205 (.a(w1133), .b(w204), .x(w649) );
	dmg_nand g1206 (.a(w188), .b(w508), .x(w1184) );
	dmg_nand g1207 (.a(w42), .b(w188), .x(w336) );
	dmg_nor3 g1208 (.a(w1025), .b(w991), .c(w990), .x(w1026) );
	dmg_nor3 g1209 (.a(w1025), .b(w980), .c(w990), .x(w992) );
	dmg_nor3 g1210 (.a(w1025), .b(w1024), .c(w979), .x(w1028) );
	dmg_nor3 g1211 (.a(w1123), .b(w1024), .c(w990), .x(w221) );
	dmg_nor3 g1212 (.a(w1123), .b(w980), .c(w979), .x(w274) );
	dmg_nor3 g1213 (.a(w1123), .b(w980), .c(w990), .x(w989) );
	dmg_nor3 g1214 (.a(w75), .b(w1016), .c(w77), .x(w78) );
	dmg_nor3 g1215 (.a(w1123), .b(w1024), .c(w979), .x(w849) );
	dmg_nor3 g1216 (.a(w70), .b(w27), .c(w163), .x(w164) );
	dmg_nor3 g1217 (.a(w766), .b(w1016), .c(w510), .x(w1187) );
	dmg_nor3 g1218 (.a(w955), .b(w70), .c(w27), .x(w26) );
	dmg_nor3 g1219 (.a(w24), .b(w1016), .c(w1112), .x(w1307) );
	dmg_nor3 g1220 (.a(w1025), .b(w980), .c(w979), .x(w978) );
	dmg_nor3 g1221 (.a(w72), .b(w70), .c(w342), .x(w73) );
	dmg_nor3 g1222 (.a(w1129), .b(w1130), .c(w1194), .x(w985) );
	dmg_nor3 g1223 (.a(w500), .b(w1016), .c(w502), .x(w1295) );
	dmg_nor3 g1224 (.a(w1299), .b(w1298), .c(w432), .x(w431) );
	dmg_nor3 g1225 (.a(w1233), .b(w70), .c(w348), .x(w543) );
	dmg_nor3 g1226 (.a(w734), .b(w1271), .c(w1270), .x(w687) );
	dmg_nor3 g1227 (.a(w70), .b(w349), .c(w676), .x(w677) );
	dmg_nor3 g1228 (.a(w70), .b(w348), .c(w603), .x(w602) );
	dmg_nor3 g1229 (.a(w70), .b(w348), .c(w661), .x(w662) );
	dmg_nand_latch g1230 (.nr(w324), .ns(w892), .nq(w325) );
	dmg_nand g1231 (.a(w188), .b(w1232), .x(w322) );
	dmg_not g1232 (.a(w306), .x(w1327) );
	dmg_dffsr g1233 (.nset1(w1323), .nset2(w1323), .d(w1097), .q(w306), .nres(w1322), .clk(w1042) );
	dmg_not6 g1234 (.a(w114), .x(w44) );
	dmg_nor3 g1235 (.a(w1171), .b(w416), .c(w922), .x(w1181) );
	dmg_fa g1236 (.cin(w425), .s(w794), .cout(w424), .a(w470), .b(w793) );
	dmg_fa g1237 (.cin(w424), .s(w890), .cout(w423), .a(w252), .b(w253) );
	dmg_fa g1238 (.cin(w231), .s(w418), .cout(w813), .a(w942), .b(w814) );
	dmg_fa g1239 (.cin(w776), .s(w775), .cout(w1401), .a(w772), .b(w773) );
	dmg_fa g1240 (.cin(w1229), .s(w1141), .cout(w1011), .a(w937), .b(w936) );
	dmg_fa g1241 (.cin(w1401), .s(w1230), .cout(w1229), .a(w1039), .b(w879) );
	dmg_fa g1242 (.cin(w813), .s(w812), .cout(w425), .a(w426), .b(w802) );
	dmg_fa g1243 (.cin(w423), .s(w422), .cout(w776), .a(w777), .b(w1403) );
	dmg_fa g1244 (.cin(w1198), .s(w1041), .cout(w1040), .a(w874), .b(w873) );
	dmg_fa g1245 (.cin(w1011), .s(w1012), .cout(w1198), .a(w934), .b(w935) );
	dmg_fa g1246 (.cin(w1040), .s(w1097), .cout(w1098), .a(w1400), .b(w1399) );
	dmg_aon222 g1247 (.a0(w527), .a1(w528), .b0(w724), .b1(w655), .c0(w654), .c1(w593), .x(w653) );
	dmg_aon222 g1248 (.a0(w724), .a1(w528), .b0(w654), .b1(w655), .c0(w592), .c1(w593), .x(w722) );
	dmg_aon22 g1249 (.a0(w134), .a1(w135), .b0(w135), .b1(w622), .x(w623) );
	dmg_aon222222 g1250 (.a0(w850), .a1(w849), .b0(w220), .b1(w221), .c0(w278), .c1(w978), .d0(w1017), .d1(w992), .e0(w277), .e1(w1028), .f0(w1030), .f1(w1026), .x(w1076) );
	dmg_aon2222 g1251 (.a0(w275), .a1(w274), .b0(w273), .b1(w989), .c0(w848), .c1(w849), .d0(w222), .d1(w221), .x(w1079) );
	dmg_aon2222 g1252 (.a0(w1063), .a1(w978), .b0(w993), .b1(w992), .c0(w1023), .c1(w1028), .d0(w1027), .d1(w1026), .x(w1078) );
	dmg_aon2222 g1253 (.a0(w633), .a1(w634), .b0(w497), .b1(w1315), .c0(w491), .c1(w490), .d0(w1313), .d1(w1314), .x(w1306) );
	dmg_aon2222 g1254 (.a0(w903), .a1(w33), .b0(w32), .b1(w1305), .c0(w896), .c1(w895), .d0(w900), .d1(w901), .x(w41) );
	dmg_notif1 g1255 (.ena(w587), .a(w577), .x(w180) );
	dmg_notif1 g1256 (.ena(w587), .a(w762), .x(w187) );
	dmg_notif1 g1257 (.ena(w587), .a(w763), .x(w229) );
	dmg_notif1 g1258 (.ena(w587), .a(w1167), .x(w29) );
	dmg_notif1 g1259 (.ena(w587), .a(w1168), .x(w16) );
	dmg_notif1 g1260 (.ena(w587), .a(w379), .x(w333) );
	dmg_notif1 g1261 (.ena(w587), .a(w517), .x(w183) );
	dmg_notif1 g1262 (.ena(w587), .a(w651), .x(w55) );
	dmg_not g1263 (.a(w144), .x(w779) );
	dmg_notif1 g1264 (.ena(w116), .a(w439), .x(w333) );
	dmg_nand5 g1265 (.a(w134), .b(w133), .c(w129), .d(w1071), .e(w841), .x(w840) );
	dmg_nand5 g1266 (.a(w964), .b(w583), .c(w112), .d(w807), .e(w808), .x(w1211) );
	dmg_nand5 g1267 (.a(w506), .b(w355), .c(w91), .d(w357), .e(w1222), .x(w92) );
	dmg_nand5 g1268 (.a(w442), .b(w443), .c(w156), .d(w545), .e(w474), .x(w473) );
	dmg_not g1269 (.a(w180), .x(w551) );
	dmg_not g1270 (.a(w1310), .x(w1309) );
	dmg_const g1271 (.q0(w20) );
	dmg_xor g1272 (.a(w231), .b(w1009), .x(w1144) );
	dmg_xor g1273 (.a(w231), .b(w307), .x(w1010) );
	dmg_xor g1274 (.a(w231), .b(w302), .x(w301) );
	dmg_xor g1275 (.a(w231), .b(w1088), .x(w875) );
	dmg_xor g1276 (.a(w231), .b(w269), .x(w268) );
	dmg_xor g1277 (.a(w231), .b(w800), .x(w870) );
	dmg_xor g1278 (.a(w231), .b(w869), .x(w866) );
	dmg_xor g1279 (.a(w231), .b(w266), .x(w943) );
	dmg_xor g1280 (.a(w231), .b(w801), .x(w267) );
	dmg_xor g1281 (.a(w231), .b(w878), .x(w419) );
	dmg_and3 g1282 (.a(w1094), .b(w1093), .c(w1031), .x(w1032) );
	dmg_and3 g1283 (.a(w289), .b(w291), .c(w290), .x(w309) );
	dmg_and3 g1284 (.a(w949), .b(w310), .c(w1086), .x(w1145) );
	dmg_and3 g1285 (.a(w293), .b(w1324), .c(w1101), .x(w1042) );
	dmg_and3 g1286 (.a(w1224), .b(w729), .c(w457), .x(w560) );
	dmg_and3 g1287 (.a(w374), .b(w375), .c(w1248), .x(w1243) );
	dmg_xor g1288 (.a(w231), .b(w232), .x(w882) );
	dmg_and3 g1289 (.a(w611), .b(w738), .c(w682), .x(w683) );
	dmg_and g1290 (.a(w911), .b(w188), .x(w656) );
	dmg_and g1291 (.a(w941), .b(w940), .x(w1364) );
	dmg_and g1292 (.a(w293), .b(w1324), .x(w1100) );
	dmg_not4 g1293 (.a(w140), .x(w141) );
	dmg_and3 g1294 (.a(w1382), .b(w335), .c(w1383), .x(w1389) );
	dmg_xnor g1295 (.x(w1390), .a(w481), .b(w482) );
	dmg_nand3 g1296 (.a(w1102), .b(w1092), .c(w948), .x(w1101) );
	dmg_or4 g1297 (.a(w111), .b(w717), .c(w112), .d(w672), .x(w1209) );
	dmg_or4 g1298 (.a(w716), .b(w583), .c(w112), .d(w672), .x(w671) );
	dmg_or4 g1299 (.a(w787), .b(w788), .c(w785), .d(w784), .x(w886) );
	dmg_nor5 g1300 (.a(w134), .b(w1283), .c(w341), .d(w484), .e(w485), .x(w843) );
	dmg_nor5 g1301 (.a(w134), .b(w133), .c(w129), .d(w1071), .e(w841), .x(w620) );
	dmg_nor5 g1302 (.a(w506), .b(w355), .c(w91), .d(w357), .e(w1222), .x(w1220) );
	dmg_nor5 g1303 (.a(w506), .b(w354), .c(w353), .d(w350), .e(w363), .x(w761) );
	dmg_and4 g1304 (.a(w208), .b(w316), .c(w63), .d(w209), .x(w320) );
	dmg_and4 g1305 (.a(w208), .b(w317), .c(w63), .d(w209), .x(w318) );
	dmg_or3 g1306 (.a(w579), .b(w587), .c(w586), .x(w710) );
	dmg_dffrnq_comp g1307 (.nr2(w40), .nr1(w40), .d(w898), .ck(w39), .cck(w650), .q(w899), .nq(w898) );
	dmg_dffrnq_comp g1308 (.nr2(w40), .nr1(w40), .d(w897), .ck(w898), .cck(w899), .q(w896), .nq(w897) );
	dmg_dffrnq_comp g1309 (.nr2(w632), .nr1(w632), .d(w493), .ck(w494), .cck(w495), .q(w492), .nq(w493) );
	dmg_dffrnq_comp g1310 (.nr2(w632), .nr1(w632), .d(w1312), .ck(w493), .cck(w492), .q(w491), .nq(w1312) );
	dmg_not g1311 (.a(w495), .x(w496) );
	dmg_or3 g1312 (.a(w70), .b(w511), .c(w761), .x(w931) );
	dmg_or3 g1313 (.a(w70), .b(w1207), .c(w410), .x(w409) );
	dmg_or3 g1314 (.a(w685), .b(w687), .c(w688), .x(w679) );
	dmg_or3 g1315 (.a(w371), .b(w431), .c(w430), .x(w437) );
	dmg_or3 g1316 (.a(w816), .b(w985), .c(w986), .x(w135) );
	dmg_or3 g1317 (.a(w70), .b(w1080), .c(w843), .x(w844) );
	dmg_not g1318 (.a(w570), .x(w237) );
	dmg_nor4 g1319 (.a(w863), .b(w985), .c(w342), .d(w70), .x(w343) );
	dmg_nor4 g1320 (.a(w1394), .b(w431), .c(w27), .d(w70), .x(w885) );
	dmg_not g1321 (.a(w371), .x(w370) );
	dmg_nor5 g1322 (.a(w442), .b(w443), .c(w156), .d(w545), .e(w474), .x(w778) );
	dmg_nor5 g1323 (.a(w442), .b(w441), .c(w214), .d(w855), .e(w534), .x(w533) );
	dmg_or g1324 (.a(w829), .b(w44), .x(w487) );
	dmg_nor4 g1325 (.a(w678), .b(w687), .c(w349), .d(w70), .x(w684) );
	dmg_and3 g1326 (.a(w1003), .b(w1004), .c(w1043), .x(w344) );
	dmg_nor6 g1327 (.a(w672), .b(w111), .c(w110), .d(w104), .e(w103), .f(w673), .x(w1356) );
	dmg_or4 g1328 (.a(w21), .b(w70), .c(w22), .d(w533), .x(w1317) );
	dmg_and4 g1329 (.a(w808), .b(w114), .c(w113), .d(w959), .x(w115) );
endmodule // APU