module APU (  cclk, clk2, clk4, clk6, clk7, clk9, n_reset2, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], cpu_wakeup, n_DRV_HIGH_a[7], n_INPUT_a[7], DRV_LOW_a[7], n_DRV_HIGH_a[6], n_INPUT_a[6], DRV_LOW_a[6], n_DRV_HIGH_a[5], n_INPUT_a[5], DRV_LOW_a[5], n_DRV_HIGH_a[4], n_INPUT_a[4], DRV_LOW_a[4], n_DRV_HIGH_a[3], n_INPUT_a[3], DRV_LOW_a[3], n_DRV_HIGH_a[2], n_INPUT_a[2], DRV_LOW_a[2], n_DRV_HIGH_a[1], n_INPUT_a[1], DRV_LOW_a[1], n_DRV_HIGH_a[0], n_INPUT_a[0], DRV_LOW_a[0], n_sout_topad, n_DRV_HIGH_sin, n_ENA_PU_sin, DRV_LOW_sin, n_DRV_HIGH_sck, sck_dir, DRV_LOW_sck, n_DRV_HIGH_p10, CONST0, n_p10, DRV_LOW_p10, n_DRV_HIGH_p11, n_p11, DRV_LOW_p11, n_DRV_HIGH_p12, n_p12, DRV_LOW_p12, n_DRV_HIGH_p13, n_p13, DRV_LOW_p13, n_DRV_HIGH_p14, DRV_LOW_p14, n_DRV_HIGH_p15, DRV_LOW_p15, dma_a[0], dma_a[4], dma_a[2], dma_a[6], dma_a[1], dma_a[5], dma_a[3], dma_a[7], soc_wr, soc_rd, lfo_512Hz, ser_out, serial_tick, test_1, test_2, n_ext_addr_en, ch3_active, wave_a[2], wave_a[3], wave_a[0], wave_a[1], wave_rd[0], wave_rd[1], wave_rd[2], wave_rd[3], wave_rd[4], wave_rd[5], wave_rd[6], wave_rd[7], n_wave_wr, wave_bl_pch, n_wave_rd, addr_latch, int_jp, FF60_D1, ffxx, n_ch1_amp_en, n_ch2_amp_en, n_ch3_amp_en, n_ch4_amp_en, ch1_out[0], ch1_out[1], ch1_out[2], ch1_out[3], ch2_out[0], ch2_out[1], ch2_out[2], ch2_out[3], ch3_out[0], ch3_out[1], ch3_out[2], ch3_out[3], ch4_out[0], ch4_out[1], ch4_out[2], ch4_out[3], r_vin_en, rmixer[0], rmixer[1], rmixer[2], rmixer[3], l_vin_en, lmixer[0], lmixer[1], lmixer[2], lmixer[3], n_rvolume[2], n_rvolume[1], n_rvolume[0], n_lvolume[2], n_lvolume[1], n_lvolume[0], from_mmio_unk1);

	input wire cclk;
	input wire clk2;
	input wire clk4;
	input wire clk6;
	input wire clk7;
	input wire clk9;
	input wire n_reset2;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	output wire cpu_wakeup;
	output wire n_DRV_HIGH_a[7];
	input wire n_INPUT_a[7];
	output wire DRV_LOW_a[7];
	output wire n_DRV_HIGH_a[6];
	input wire n_INPUT_a[6];
	output wire DRV_LOW_a[6];
	output wire n_DRV_HIGH_a[5];
	input wire n_INPUT_a[5];
	output wire DRV_LOW_a[5];
	output wire n_DRV_HIGH_a[4];
	input wire n_INPUT_a[4];
	output wire DRV_LOW_a[4];
	output wire n_DRV_HIGH_a[3];
	input wire n_INPUT_a[3];
	output wire DRV_LOW_a[3];
	output wire n_DRV_HIGH_a[2];
	input wire n_INPUT_a[2];
	output wire DRV_LOW_a[2];
	output wire n_DRV_HIGH_a[1];
	input wire n_INPUT_a[1];
	output wire DRV_LOW_a[1];
	output wire n_DRV_HIGH_a[0];
	input wire n_INPUT_a[0];
	output wire DRV_LOW_a[0];
	output wire n_sout_topad;
	output wire n_DRV_HIGH_sin;
	output wire n_ENA_PU_sin;
	output wire DRV_LOW_sin;
	output wire n_DRV_HIGH_sck;
	input wire sck_dir;
	output wire DRV_LOW_sck;
	output wire n_DRV_HIGH_p10;
	input wire CONST0;
	input wire n_p10;
	output wire DRV_LOW_p10;
	output wire n_DRV_HIGH_p11;
	input wire n_p11;
	output wire DRV_LOW_p11;
	output wire n_DRV_HIGH_p12;
	input wire n_p12;
	output wire DRV_LOW_p12;
	output wire n_DRV_HIGH_p13;
	input wire n_p13;
	output wire DRV_LOW_p13;
	output wire n_DRV_HIGH_p14;
	output wire DRV_LOW_p14;
	output wire n_DRV_HIGH_p15;
	output wire DRV_LOW_p15;
	input wire dma_a[0];
	input wire dma_a[4];
	input wire dma_a[2];
	input wire dma_a[6];
	input wire dma_a[1];
	input wire dma_a[5];
	input wire dma_a[3];
	input wire dma_a[7];
	input wire soc_wr;
	input wire soc_rd;
	input wire lfo_512Hz;
	input wire ser_out;
	input wire serial_tick;
	input wire test_1;
	input wire test_2;
	input wire n_ext_addr_en;
	output wire ch3_active;
	output wire wave_a[2];
	output wire wave_a[3];
	output wire wave_a[0];
	output wire wave_a[1];
	input wire wave_rd[0];
	input wire wave_rd[1];
	input wire wave_rd[2];
	input wire wave_rd[3];
	input wire wave_rd[4];
	input wire wave_rd[5];
	input wire wave_rd[6];
	input wire wave_rd[7];
	output wire n_wave_wr;
	output wire wave_bl_pch;
	output wire n_wave_rd;
	input wire addr_latch;
	output wire int_jp;
	output wire FF60_D1;
	input wire ffxx;
	output wire n_ch1_amp_en;
	output wire n_ch2_amp_en;
	output wire n_ch3_amp_en;
	output wire n_ch4_amp_en;
	output wire ch1_out[0];
	output wire ch1_out[1];
	output wire ch1_out[2];
	output wire ch1_out[3];
	output wire ch2_out[0];
	output wire ch2_out[1];
	output wire ch2_out[2];
	output wire ch2_out[3];
	output wire ch3_out[0];
	output wire ch3_out[1];
	output wire ch3_out[2];
	output wire ch3_out[3];
	output wire ch4_out[0];
	output wire ch4_out[1];
	output wire ch4_out[2];
	output wire ch4_out[3];
	output wire r_vin_en;
	output wire rmixer[0];
	output wire rmixer[1];
	output wire rmixer[2];
	output wire rmixer[3];
	output wire l_vin_en;
	output wire lmixer[0];
	output wire lmixer[1];
	output wire lmixer[2];
	output wire lmixer[3];
	output wire n_rvolume[2];
	output wire n_rvolume[1];
	output wire n_rvolume[0];
	output wire n_lvolume[2];
	output wire n_lvolume[1];
	output wire n_lvolume[0];
	input wire from_mmio_unk1;

endmodule // APU