module OAM (  n_oamb[0], n_oamb[1], n_oamb[2], n_oamb[3], n_oamb[4], n_oamb[5], n_oamb[6], n_oamb[7], oam_bl_pch, oa[1], oa[2], oa[3], oa[4], oa[5], oa[6], oa[7], n_oam_rd, n_oamb_wr, n_oama_wr, n_oama[0], n_oama[1], n_oama[2], n_oama[3], n_oama[4], n_oama[5], n_oama[6], n_oama[7]);

	inout wire n_oamb[0];
	inout wire n_oamb[1];
	inout wire n_oamb[2];
	inout wire n_oamb[3];
	inout wire n_oamb[4];
	inout wire n_oamb[5];
	inout wire n_oamb[6];
	inout wire n_oamb[7];
	input wire oam_bl_pch;
	input wire oa[1];
	input wire oa[2];
	input wire oa[3];
	input wire oa[4];
	input wire oa[5];
	input wire oa[6];
	input wire oa[7];
	input wire n_oam_rd;
	input wire n_oamb_wr;
	input wire n_oama_wr;
	inout wire n_oama[0];
	inout wire n_oama[1];
	inout wire n_oama[2];
	inout wire n_oama[3];
	inout wire n_oama[4];
	inout wire n_oama[5];
	inout wire n_oama[6];
	inout wire n_oama[7];

endmodule // OAM