module dmgcpu (  sck, md, d, p13, p12, p11, p10, sin, n_res, t2, t1, a, n_cs, n_rd, n_wr, phi, ck1, ck2, sout, p14, p15, so2, so1, s, fr, cpl, st, cp, cpg, ld0, ld1, n_mwr, ma, n_mrd, n_mcs, vin);

	inout wire sck;
	inout wire [7:0] md;
	inout wire [7:0] d;
	inout wire p13;
	inout wire p12;
	inout wire p11;
	inout wire p10;
	inout wire sin;
	input wire n_res;
	input wire t2;
	input wire t1;
	inout wire [15:0] a;
	output wire n_cs;
	inout wire n_rd;
	inout wire n_wr;
	output wire phi;
	input wire ck1;
	output wire ck2;
	output wire sout;
	output wire p14;
	output wire p15;
	output wire so2;
	output wire so1;
	output wire s;
	output wire fr;
	output wire cpl;
	output wire st;
	output wire cp;
	output wire cpg;
	output wire ld0;
	output wire ld1;
	inout wire n_mwr;
	output wire [12:0] ma;
	inout wire n_mrd;
	inout wire n_mcs;
	input wire vin;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;

	assign sck = w1;
	assign md[0] = w2;
	assign md[1] = w3;
	assign md[2] = w4;
	assign md[3] = w5;
	assign md[4] = w6;
	assign md[5] = w7;
	assign md[6] = w8;
	assign md[7] = w9;
	assign d[7] = w10;
	assign d[6] = w11;
	assign d[5] = w12;
	assign d[4] = w13;
	assign d[3] = w14;
	assign d[2] = w15;
	assign d[1] = w16;
	assign d[0] = w17;
	assign p13 = w18;
	assign p12 = w19;
	assign p11 = w20;
	assign p10 = w21;
	assign sin = w22;
	assign w23 = n_res;
	assign w24 = t2;
	assign w25 = t1;
	assign a[15] = w26;
	assign a[14] = w27;
	assign a[13] = w28;
	assign a[12] = w29;
	assign a[11] = w30;
	assign a[10] = w31;
	assign a[9] = w32;
	assign a[8] = w33;
	assign a[7] = w34;
	assign a[6] = w35;
	assign a[5] = w36;
	assign a[4] = w37;
	assign a[3] = w38;
	assign a[2] = w39;
	assign a[1] = w40;
	assign a[0] = w41;
	assign n_cs = w42;
	assign n_rd = w43;
	assign n_wr = w44;
	assign phi = w45;
	assign w46 = ck1;
	assign ck2 = w47;
	assign sout = w48;
	assign p14 = w49;
	assign p15 = w50;
	assign so2 = w51;
	assign so1 = w52;
	assign s = w53;
	assign fr = w54;
	assign cpl = w55;
	assign st = w56;
	assign cp = w57;
	assign cpg = w58;
	assign ld0 = w59;
	assign ld1 = w60;
	assign n_mwr = w61;
	assign ma[8] = w62;
	assign ma[9] = w63;
	assign ma[11] = w64;
	assign n_mrd = w65;
	assign ma[10] = w66;
	assign n_mcs = w67;
	assign ma[12] = w68;
	assign ma[7] = w69;
	assign ma[6] = w70;
	assign ma[5] = w71;
	assign ma[4] = w72;
	assign ma[3] = w73;
	assign ma[2] = w74;
	assign ma[1] = w75;
	assign ma[0] = w76;
	assign w77 = vin;

	// Instances

	dmgcpu_IOBUF_B pad_d6 (.DRV_LOW(w318), .n_INPUT(w317), .n_ENA_PU(w315), .n_DRV_HIGH(w316), .PAD_IO(w11) );
	dmgcpu_IOBUF_B pad_d7 (.DRV_LOW(w314), .n_INPUT(w313), .n_ENA_PU(w315), .n_DRV_HIGH(w312), .PAD_IO(w10) );
	dmgcpu_IOBUF_B pad_md7 (.DRV_LOW(w289), .n_INPUT(w288), .n_ENA_PU(w290), .n_DRV_HIGH(w287), .PAD_IO(w9) );
	dmgcpu_IOBUF_B pad_md6 (.DRV_LOW(w293), .n_INPUT(w292), .n_ENA_PU(w290), .n_DRV_HIGH(w291), .PAD_IO(w8) );
	dmgcpu_IOBUF_B pad_md5 (.DRV_LOW(w296), .n_INPUT(w295), .n_ENA_PU(w290), .n_DRV_HIGH(w294), .PAD_IO(w7) );
	dmgcpu_IOBUF_B pad_md4 (.DRV_LOW(w299), .n_INPUT(w298), .n_ENA_PU(w290), .n_DRV_HIGH(w297), .PAD_IO(w6) );
	dmgcpu_IOBUF_B pad_md3 (.DRV_LOW(w302), .n_INPUT(w301), .n_ENA_PU(w290), .n_DRV_HIGH(w300), .PAD_IO(w5) );
	dmgcpu_IOBUF_B pad_md2 (.DRV_LOW(w305), .n_INPUT(w304), .n_ENA_PU(w290), .n_DRV_HIGH(w303), .PAD_IO(w4) );
	dmgcpu_IOBUF_B pad_md1 (.DRV_LOW(w308), .n_INPUT(w307), .n_ENA_PU(w290), .n_DRV_HIGH(w306), .PAD_IO(w3) );
	dmgcpu_IOBUF_B pad_md0 (.DRV_LOW(w310), .n_INPUT(w311), .n_ENA_PU(w290), .n_DRV_HIGH(w309), .PAD_IO(w2) );
	dmgcpu_IOBUF_C pad_sck (.n_DRV_HIGH(w254), .n_ENA_PU(w255), .DRV_LOW(w257), .n_INPUT(w256), .PAD_IO(w1) );
	dmgcpu_IOBUF_B pad_d5 (.PAD_IO(w12), .DRV_LOW(w321), .n_DRV_HIGH(w319), .n_ENA_PU(w315), .n_INPUT(w320) );
	dmgcpu_IOBUF_B pad_d4 (.PAD_IO(w13), .DRV_LOW(w324), .n_DRV_HIGH(w322), .n_ENA_PU(w315), .n_INPUT(w323) );
	dmgcpu_IOBUF_B pad_d3 (.PAD_IO(w14), .DRV_LOW(w327), .n_DRV_HIGH(w325), .n_ENA_PU(w315), .n_INPUT(w326) );
	dmgcpu_IOBUF_B pad_d2 (.PAD_IO(w15), .DRV_LOW(w330), .n_DRV_HIGH(w328), .n_ENA_PU(w315), .n_INPUT(w329) );
	dmgcpu_IOBUF_B pad_d1 (.PAD_IO(w16), .DRV_LOW(w333), .n_DRV_HIGH(w331), .n_ENA_PU(w315), .n_INPUT(w332) );
	dmgcpu_IOBUF_B pad_d0 (.PAD_IO(w17), .n_DRV_HIGH(w334), .n_ENA_PU(w315), .n_INPUT(w335) );
	dmgcpu_IOBUF_B pad_sin (.PAD_IO(w22), .DRV_LOW(w253), .n_ENA_PU(w251), .n_DRV_HIGH(w250), .n_INPUT(w252) );
	dmgcpu_IOBUF_B pad_p10 (.PAD_IO(w21), .DRV_LOW(w261), .n_ENA_PU(w259), .n_DRV_HIGH(w258), .n_INPUT(w260) );
	dmgcpu_IOBUF_B pad_p11 (.PAD_IO(w20), .DRV_LOW(w264), .n_ENA_PU(w259), .n_DRV_HIGH(w262), .n_INPUT(w263) );
	dmgcpu_IOBUF_B pad_p12 (.PAD_IO(w19), .DRV_LOW(w267), .n_ENA_PU(w259), .n_DRV_HIGH(w265), .n_INPUT(w266) );
	dmgcpu_IOBUF_B pad_p13 (.PAD_IO(w18), .DRV_LOW(w270), .n_ENA_PU(w259), .n_DRV_HIGH(w268), .n_INPUT(w269) );
	dmgcpu_IBUF_A pad_t1 (.n_INPUT(w247), .PAD_IN(w25) );
	dmgcpu_IBUF_A pad_t2 (.n_INPUT(w248), .PAD_IN(w24) );
	dmgcpu_IBUF_A pad_nres (.n_INPUT(w79), .PAD_IN(w23) );
	dmgcpu_IOBUF_A pad_a15 (.PAD_IO(w26), .n_DRV_HIGH(w192), .DRV_LOW(w194), .n_INPUT(w193) );
	dmgcpu_IOBUF_A pad_a14 (.PAD_IO(w27), .n_DRV_HIGH(w195), .DRV_LOW(w197), .n_INPUT(w196) );
	dmgcpu_IOBUF_A pad_a13 (.PAD_IO(w28), .n_DRV_HIGH(w198), .DRV_LOW(w200), .n_INPUT(w199) );
	dmgcpu_IOBUF_A pad_a12 (.PAD_IO(w29), .n_DRV_HIGH(w201), .DRV_LOW(w203), .n_INPUT(w202) );
	dmgcpu_IOBUF_A pad_a11 (.PAD_IO(w30), .n_DRV_HIGH(w204), .DRV_LOW(w206), .n_INPUT(w205) );
	dmgcpu_IOBUF_A pad_a10 (.PAD_IO(w31), .n_DRV_HIGH(w207), .DRV_LOW(w209), .n_INPUT(w208) );
	dmgcpu_IOBUF_A pad_a9 (.PAD_IO(w32), .n_DRV_HIGH(w210), .DRV_LOW(w212), .n_INPUT(w211) );
	dmgcpu_IOBUF_A pad_a8 (.PAD_IO(w33), .n_DRV_HIGH(w213), .DRV_LOW(w215), .n_INPUT(w214) );
	dmgcpu_IOBUF_A pad_a7 (.PAD_IO(w34), .n_DRV_HIGH(w216), .DRV_LOW(w218), .n_INPUT(w217) );
	dmgcpu_IOBUF_A pad_a6 (.PAD_IO(w35), .n_DRV_HIGH(w219), .DRV_LOW(w221), .n_INPUT(w220) );
	dmgcpu_IOBUF_A pad_a5 (.PAD_IO(w36), .n_DRV_HIGH(w222), .DRV_LOW(w224), .n_INPUT(w223) );
	dmgcpu_IOBUF_A pad_a4 (.PAD_IO(w37), .n_DRV_HIGH(w225), .DRV_LOW(w227), .n_INPUT(w226) );
	dmgcpu_IOBUF_A pad_a3 (.PAD_IO(w38), .n_DRV_HIGH(w228), .DRV_LOW(w230), .n_INPUT(w229) );
	dmgcpu_IOBUF_A pad_a2 (.PAD_IO(w39), .n_DRV_HIGH(w231), .DRV_LOW(w233), .n_INPUT(w232) );
	dmgcpu_IOBUF_A pad_a1 (.PAD_IO(w40), .n_DRV_HIGH(w234), .DRV_LOW(w236), .n_INPUT(w235) );
	dmgcpu_IOBUF_A pad_a0 (.PAD_IO(w41), .n_DRV_HIGH(w237), .DRV_LOW(w239), .n_INPUT(w238) );
	dmgcpu_IOBUF_A pad_nrd (.PAD_IO(w43), .n_DRV_HIGH(w241), .DRV_LOW(w243), .n_INPUT(w242) );
	dmgcpu_IOBUF_A pad_nwr (.PAD_IO(w44), .n_DRV_HIGH(w244), .DRV_LOW(w246), .n_INPUT(w245) );
	dmgcpu_IOBUF_A pad_nmcs (.PAD_IO(w67), .n_DRV_HIGH(w284), .n_INPUT(w285) );
	dmgcpu_IOBUF_A pad_nmrd (.PAD_IO(w65), .DRV_LOW(w283), .n_DRV_HIGH(w281), .n_INPUT(w282) );
	dmgcpu_IOBUF_A pad_nmwr (.PAD_IO(w61), .DRV_LOW(w280), .n_DRV_HIGH(w278), .n_INPUT(w279) );
	dmgcpu_OBUF_A pad_s (.n_OUTPUT(w164), .PAD_OUT(w53) );
	dmgcpu_OBUF_A pad_fr (.n_OUTPUT(w163), .PAD_OUT(w54) );
	dmgcpu_OBUF_A pad_cpl (.n_OUTPUT(w162), .PAD_OUT(w55) );
	dmgcpu_OBUF_A pad_st (.n_OUTPUT(w161), .PAD_OUT(w56) );
	dmgcpu_OBUF_A pad_cp (.n_OUTPUT(w160), .PAD_OUT(w57) );
	dmgcpu_OBUF_A pad_cpg (.n_OUTPUT(w159), .PAD_OUT(w58) );
	dmgcpu_OBUF_A pad_m1 (.n_OUTPUT(w100) );
	dmgcpu_OBUF_A pad_ld0 (.n_OUTPUT(w158), .PAD_OUT(w59) );
	dmgcpu_OBUF_A pad_ld1 (.n_OUTPUT(w157), .PAD_OUT(w60) );
	dmgcpu_OBUF_A pad_ma8 (.n_OUTPUT(w147), .PAD_OUT(w62) );
	dmgcpu_OBUF_A pad_ma9 (.n_OUTPUT(w148), .PAD_OUT(w63) );
	dmgcpu_OBUF_A pad_ma11 (.n_OUTPUT(w146), .PAD_OUT(w64) );
	dmgcpu_OBUF_A pad_ma10 (.n_OUTPUT(w145), .PAD_OUT(w66) );
	dmgcpu_OBUF_A pad_ma12 (.n_OUTPUT(w144), .PAD_OUT(w68) );
	dmgcpu_OBUF_A pad_ma7 (.n_OUTPUT(w151), .PAD_OUT(w69) );
	dmgcpu_OBUF_A pad_ma6 (.n_OUTPUT(w149), .PAD_OUT(w70) );
	dmgcpu_OBUF_A pad_ma5 (.n_OUTPUT(w150), .PAD_OUT(w71) );
	dmgcpu_OBUF_A pad_ma4 (.n_OUTPUT(w154), .PAD_OUT(w72) );
	dmgcpu_OBUF_A pad_ma3 (.n_OUTPUT(w152), .PAD_OUT(w73) );
	dmgcpu_OBUF_A pad_ma2 (.n_OUTPUT(w153), .PAD_OUT(w74) );
	dmgcpu_OBUF_A pad_ma1 (.n_OUTPUT(w155), .PAD_OUT(w75) );
	dmgcpu_OBUF_A pad_ma0 (.n_OUTPUT(w156), .PAD_OUT(w76) );
	dmgcpu_AOBUFFER pad_so1 (.VOUT(w277), .PAD_OUT(w52) );
	dmgcpu_AOBUFFER pad_so2 (.VOUT(w276), .PAD_OUT(w51) );
	dmgcpu_OBUF_B pad_p15 (.n_DRV_HIGH(w273), .DRV_LOW(w274), .PAD_OUT(w50) );
	dmgcpu_OBUF_B pad_p14 (.DRV_LOW(w272), .n_DRV_HIGH(w271), .PAD_OUT(w49) );
	dmgcpu_IBUF_B pad_nnmi (.n_INPUT(w98) );
	dmgcpu_OBUF_A pad_ncs (.PAD_OUT(w42), .n_OUTPUT(w240) );
	dmgcpu_OBUF_A pad_phi (.PAD_OUT(w45), .n_OUTPUT(w84) );
	dmgcpu_OSC ck1_ck2 (.ENA(w87), .n_CLK(w78), .CK_IN(w46), .CK_OUT(w47) );
	dmgcpu_OBUF_A pad_sout (.PAD_OUT(w48), .n_OUTPUT(w249) );
	dmgcpu_AIBUFFER pad_vin (.VIN(w275), .PAD_IN(w77) );
	dmgcpu_PPU1 ppu1 (.a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .a[8](w117), .a[9](w118), .a[10](w119), .a[11](w120), .a[12](w121), .n_ma[12](w144), .n_ma[10](w145), .n_ma[11](w146), .n_ma[8](w147), .n_ma[9](w148), .n_ma[6](w149), .n_ma[5](w150), .n_ma[7](w151), .n_ma[3](w152), .n_ma[2](w153), .n_ma[4](w154), .n_ma[1](w155), .n_ma[0](w156), .lcd_ld1(w157), .lcd_ld0(w158), .lcd_cpg(w159), .lcd_cp(w160), .lcd_st(w161), .lcd_cpl(w162), .lcd_fr(w163), .lcd_s(w164), .CONST0(w259), .n_dma_phi(w337), .ppu_rd(w355), .ppu_wr(w356), .ppu_clk(w365), .vram_to_oam(w366), .ffxx(w395), .n_ppu_hard_reset(w396), .ff46(w397), .nma[9](w398), .fexx(w399), .nma[0](w400), .ff43(w401), .nma[4](w402), .nma[12](w403), .nma[6](w404), .nma[5](w405), .ff42(w406), .nma[11](w407), .nma[10](w408), .sprite_x_flip(w409), .nma[3](w410), .nma[2](w411), .sprite_x_match(w412), .bp_sel(w413) );
	dmgcpu_PPU2 ppu2 (.cclk(w80), .clk6(w89), .n_reset2(w93), .a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .n_oamb[0](w165), .n_oamb[1](w166), .n_oamb[2](w167), .n_oamb[3](w168), .n_oamb[4](w169), .n_oamb[5](w170), .n_oamb[6](w171), .n_oamb[7](w172), .oam_bl_pch(w173), .oa[1](w174), .oa[2](w175), .oa[3](w176), .oa[4](w177), .oa[5](w178), .oa[6](w179), .oa[7](w180), .n_oam_rd(w181), .n_oamb_wr(w182), .n_oama_wr(w183), .n_oama[0](w184), .n_oama[1](w185), .n_oama[2](w186), .n_oama[3](w187), .n_oama[4](w188), .n_oama[5](w189), .n_oama[6](w190), .n_oama[7](w191), .CONST0(w259), .n_dma_phi(w337), .dma_a[0](w338), .dma_a[4](w339), .dma_a[2](w340), .dma_a[6](w341), .dma_a[10](w342), .dma_a[1](w343), .dma_a[5](w344), .dma_a[11](w345), .dma_a[3](w346), .dma_a[7](w347), .dma_a[8](w348), .dma_a[12](w349), .dma_a[9](w350), .dma_run(w351), .soc_wr(w352), .soc_rd(w353), .ppu_rd(w355), .ppu_wr(w356), .ppu_clk(w365), .vram_to_oam(w366), .n_ppu_hard_reset(w396), .nma[9](w398), .fexx(w399), .nma[0](w400), .ff43(w401), .nma[4](w402), .nma[12](w403), .nma[6](w404), .nma[5](w405), .ff42(w406), .nma[11](w407), .nma[10](w408), .sprite_x_flip(w409), .nma[3](w410), .nma[2](w411), .sprite_x_match(w412), .bp_sel(w413) );
	dmgcpu_OAM oam (.n_oamb[0](w165), .n_oamb[1](w166), .n_oamb[2](w167), .n_oamb[3](w168), .n_oamb[4](w169), .n_oamb[5](w170), .n_oamb[6](w171), .n_oamb[7](w172), .oam_bl_pch(w173), .oa[1](w174), .oa[2](w175), .oa[3](w176), .oa[4](w177), .oa[5](w178), .oa[6](w179), .oa[7](w180), .n_oam_rd(w181), .n_oamb_wr(w182), .n_oama_wr(w183), .n_oama[0](w184), .n_oama[1](w185), .n_oama[2](w186), .n_oama[3](w187), .n_oama[4](w188), .n_oama[5](w189), .n_oama[6](w190), .n_oama[7](w191) );
	dmgcpu_HRAM hram (.clk7(w90), .a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4(w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .soc_wr(w352), .soc_rd(w353), .ffxx(w395) );
	dmgcpu_DAC dac (.vin_analog(w275), .so2_analog(w276), .so1_analog(w277) );
	dmgcpu_BootROM bootrom (.a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .a[8](w117), .a[9](w118), .a[10](w119), .a[11](w120), .a[12](w121), .a[13](w122), .a[14](w123), .a[15](w124) );
	dmgcpu_Ser ser (.n_reset2(w93), .d[5](w105), .d[6](w104), .d[7](w103), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .n_sin(w252), .sck_dir(w255), .n_sck(w256), .int_serial(w357), .sc_read(w358), .sb_read(w359), .sc_write(w360), .n_sb_write(w361), .lfo_16384Hz(w362), .ser_out(w363), .serial_tick(w364) );
	dmgcpu_ClkGen clkgen (.n_clk_in(w78), .reset(w79), .cclk(w80), .clk1(w81), .clk2(w82), .clk3(w83), .clk4(w84), .osc_stable(w85), .clk_ena(w86), .osc_ena(w87), .clk5(w88), .clk6(w89), .clk7(w90), .clk8(w91), .clk9(w92), .n_reset2(w93), .sync_reset(w94), .cpu_mreq(w95), .ext_cs_en(w96), .cpu_wr_sync(w97), .cpu_wr(w140), .test_1(w369), .n_test_reset(w374) );
	dmgcpu_MMIO mmio (.reset(w79), .clk2(w82), .clk4(w84), .osc_stable(w85), .clk_ena(w86), .osc_ena(w87), .clk6(w89), .clk9(w92), .n_reset2(w93), .cpu_wr_sync(w97), .cpu_m1(w99), .n_cpu_m1(w100), .a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .a[8](w117), .a[9](w118), .a[10](w119), .a[11](w120), .a[12](w121), .a[13](w122), .a[14](w123), .cpu_irq_trig[4](w128), .cpu_irq_ack[4](w129), .cpu_irq_trig[3](w130), .cpu_irq_ack[3](w131), .cpu_irq_trig[2](w132), .cpu_irq_ack[2](w133), .cpu_irq_trig[1](w134), .cpu_irq_ack[1](w135), .cpu_irq_trig[0](w136), .cpu_irq_ack[0](w137), .cpu_rd(w139), .cpu_wr(w140), .n_DRV_HIGH_a[14](w195), .n_INPUT_a[14](w196), .DRV_LOW_a[14](w197), .n_DRV_HIGH_a[13](w198), .n_INPUT_a[13](w199), .DRV_LOW_a[13](w200), .n_DRV_HIGH_a[12](w201), .n_INPUT_a[12](w202), .DRV_LOW_a[12](w203), .n_DRV_HIGH_a[11](w204), .n_INPUT_a[11](w205), .DRV_LOW_a[11](w206), .n_DRV_HIGH_a[10](w207), .n_INPUT_a[10](w208), .DRV_LOW_a[10](w209), .n_DRV_HIGH_a[9](w210), .n_INPUT_a[9](w211), .DRV_LOW_a[9](w212), .n_DRV_HIGH_a[8](w213), .n_INPUT_a[8](w214), .DRV_LOW_a[8](w215), .n_DRV_HIGH_nrd(w241), .n_INPUT_nrd(w242), .DRV_LOW_nrd(w243), .n_DRV_HIGH_nwr(w244), .n_INPUT_nwr(w245), .DRV_LOW_nwr(w246), .n_t1_frompad(w247), .n_t2_frompad(w248), .CONST0(w259), .n_ena_pu_db(w315), .n_dma_phi(w337), .dma_a[0](w338), .dma_a[4](w339), .dma_a[2](w340), .dma_a[6](w341), .dma_a[10](w342), .dma_a[1](w343), .dma_a[5](w344), .dma_a[11](w345), .dma_a[3](w346), .dma_a[7](w347), .dma_a[8](w348), .dma_a[12](w349), .dma_a[9](w350), .dma_run(w351), .soc_wr(w352), .soc_rd(w353), .lfo_512Hz(w354), .ppu_rd(w355), .ppu_wr(w356), .int_serial(w357), .sc_read(w358), .sb_read(w359), .sc_write(w360), .n_sb_write(w361), .lfo_16384Hz(w362), .ppu_clk(w365), .vram_to_oam(w366), .dma_a[15](w367), .non_vram_mreq(w368), .test_1(w369), .test_2(w370), .n_extdb_to_intdb(w371), .n_dblatch_to_intdb(w372), .n_intdb_to_extdb(w373), .n_test_reset(w374), .n_ext_addr_en(w375), .addr_latch(w392), .int_jp(w393), .FF60_D1(w394), .ffxx(w395), .n_ppu_hard_reset(w396), .ff46(w397) );
	dmgcpu_SM83Core core (.RESET(w79), .CLK1(w81), .CLK2(w82), .CLK3(w83), .CLK4(w84), .OSC_STABLE(w85), .CLK_ENA(w86), .OSC_ENA(w87), .CLK5(w88), .CLK6(w89), .CLK7(w90), .CLK8(w91), .CLK9(w92), .SYNC_RESET(w94), .CPU_MREQ(w95), .NMI(w98), .M1(w99), .A[0](w101), .A[1](w102), .D[7](w103), .D[6](w104), .D[5](w105), .D[4](w106), .D[3](w107), .D[2](w108), .D[1](w109), .D[0](w110), .A[2](w111), .A[3](w112), .A[4](w113), .A[5](w114), .A[6](w115), .A[7](w116), .A[8](w117), .A[9](w118), .A[10](w119), .A[11](w120), .A[12](w121), .A[13](w122), .A[14](w123), .A[15](w124), .CPU_IRQ_TRIG[7](1'b0), .CPU_IRQ_TRIG[6](1'b0), .CPU_IRQ_TRIG[5](1'b0), .CPU_IRQ_TRIG[4](w128), .CPU_IRQ_ACK[4](w129), .CPU_IRQ_TRIG[3](w130), .CPU_IRQ_ACK[3](w131), .CPU_IRQ_TRIG[2](w132), .CPU_IRQ_ACK[2](w133), .CPU_IRQ_TRIG[1](w134), .CPU_IRQ_ACK[1](w135), .CPU_IRQ_TRIG[0](w136), .CPU_IRQ_ACK[0](w137), .WAKE(w138), .RD(w139), .WR(w140), .MMIO_REQ(w141), .IPL_REQ(w142), .BUS_DISABLE(w369), .IPL_DISABLE(w370) );
	dmgcpu_Arbiter arb (.clk2(w82), .n_reset2(w93), .cpu_mreq(w95), .ext_cs_en(w96), .cpu_wr_sync(w97), .a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .a[8](w117), .a[9](w118), .a[10](w119), .a[11](w120), .a[12](w121), .a[13](w122), .a[14](w123), .a[15](w124), .cpu_wr(w140), .mmio_sel(w141), .boot_sel(w142), .n_DRV_HIGH_a[15](w192), .n_INPUT_a[15](w193), .DRV_LOW_a[15](w194), .n_cs_topad(w240), .CONST0(w259), .n_DRV_HIGH_nmwr(w278), .n_mwr(w279), .DRV_LOW_nmwr(w280), .n_DRV_HIGH_nmrd(w281), .n_mrd(w282), .DRV_LOW_nmrd(w283), .n_DRV_HIGH_nmcs(w284), .n_mcs(w285), .DRV_LOW_nmcs(w286), .n_DRV_HIGH_md[7](w287), .n_md_frompad[7](w288), .DRV_LOW_md[7](w289), .n_md_ena_pu(w290), .n_DRV_HIGH_md[6](w291), .n_md_frompad[6](w292), .DRV_LOW_md[6](w293), .n_DRV_HIGH_md[5](w294), .n_md_frompad[5](w295), .DRV_LOW_md[5](w296), .n_DRV_HIGH_md[4](w297), .n_md_frompad[4](w298), .DRV_LOW_md[4](w299), .n_DRV_HIGH_md[3](w300), .n_md_frompad[3](w301), .DRV_LOW_md[3](w302), .n_DRV_HIGH_md[2](w303), .n_md_frompad[2](w304), .DRV_LOW_md[2](w305), .n_DRV_HIGH_md[1](w306), .n_md_frompad[1](w307), .DRV_LOW_md[1](w308), .n_DRV_HIGH_md[0](w309), .DRV_LOW_md[0](w310), .n_md_frompad[0](w311), .n_DRV_HIGH_d[7](w312), .n_db_frompad[7](w313), .DRV_LOW_d[7](w314), .n_ena_pu_db(w315), .n_DRV_HIGH_d[6](w316), .n_db_frompad[6](w317), .DRV_LOW_d[6](w318), .n_DRV_HIGH_d[5](w319), .n_db_frompad[5](w320), .DRV_LOW_d[5](w321), .n_DRV_HIGH_d[4](w322), .n_db_frompad[4](w323), .DRV_LOW_d[4](w324), .n_DRV_HIGH_d[3](w325), .n_db_frompad[3](w326), .DRV_LOW_d[3](w327), .n_DRV_HIGH_d[2](w328), .n_db_frompad[2](w329), .DRV_LOW_d[2](w330), .n_DRV_HIGH_d[1](w331), .n_db_frompad[1](w332), .DRV_LOW_d[1](w333), .n_DRV_HIGH_d[0](w334), .n_db_frompad[0](w335), .DRV_LOW_a[0](w336), .soc_wr(w352), .soc_rd(w353), .vram_to_oam(w366), .dma_a[15](w367), .non_vram_mreq(w368), .test_1(w369), .n_extdb_to_intdb(w371), .n_dblatch_to_intdb(w372), .n_intdb_to_extdb(w373), .ffxx(w395), .n_ppu_hard_reset(w396) );
	dmgcpu_APU apu (.cclk(w80), .clk2(w82), .clk4(w84), .clk6(w89), .clk7(w90), .clk9(w92), .n_reset2(w93), .a[0](w101), .a[1](w102), .d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .a[2](w111), .a[3](w112), .a[4](w113), .a[5](w114), .a[6](w115), .a[7](w116), .cpu_wakeup(w138), .n_DRV_HIGH_a[7](w216), .n_INPUT_a[7](w217), .DRV_LOW_a[7](w218), .n_DRV_HIGH_a[6](w219), .n_INPUT_a[6](w220), .DRV_LOW_a[6](w221), .n_DRV_HIGH_a[5](w222), .n_INPUT_a[5](w223), .DRV_LOW_a[5](w224), .n_DRV_HIGH_a[4](w225), .n_INPUT_a[4](w226), .DRV_LOW_a[4](w227), .n_DRV_HIGH_a[3](w228), .n_INPUT_a[3](w229), .DRV_LOW_a[3](w230), .n_DRV_HIGH_a[2](w231), .n_INPUT_a[2](w232), .DRV_LOW_a[2](w233), .n_DRV_HIGH_a[1](w234), .n_INPUT_a[1](w235), .DRV_LOW_a[1](w236), .n_DRV_HIGH_a[0](w237), .n_INPUT_a[0](w238), .DRV_LOW_a[0](w239), .n_sout_topad(w249), .n_DRV_HIGH_sin(w250), .n_ENA_PU_sin(w251), .DRV_LOW_sin(w253), .n_DRV_HIGH_sck(w254), .sck_dir(w255), .DRV_LOW_sck(w257), .n_DRV_HIGH_p10(w258), .CONST0(w259), .n_p10(w260), .DRV_LOW_p10(w261), .n_DRV_HIGH_p11(w262), .n_p11(w263), .DRV_LOW_p11(w264), .n_DRV_HIGH_p12(w265), .n_p12(w266), .DRV_LOW_p12(w267), .n_DRV_HIGH_p13(w268), .n_p13(w269), .DRV_LOW_p13(w270), .n_DRV_HIGH_p14(w271), .DRV_LOW_p14(w272), .n_DRV_HIGH_p15(w273), .DRV_LOW_p15(w274), .dma_a[0](w338), .dma_a[4](w339), .dma_a[2](w340), .dma_a[6](w341), .dma_a[1](w343), .dma_a[5](w344), .dma_a[3](w346), .dma_a[7](w347), .soc_wr(w352), .soc_rd(w353), .lfo_512Hz(w354), .ser_out(w363), .serial_tick(w364), .test_1(w369), .test_2(w370), .n_ext_addr_en(w375), .ch3_active(w376), .wave_a[2](w377), .wave_a[3](w378), .wave_a[0](w379), .wave_a[1](w380), .wave_rd[0](w381), .wave_rd[1](w382), .wave_rd[2](w383), .wave_rd[3](w384), .wave_rd[4](w385), .wave_rd[5](w386), .wave_rd[6](w387), .wave_rd[7](w388), .n_wave_wr(w389), .wave_bl_pch(w390), .n_wave_rd(w391), .addr_latch(w392), .int_jp(w393), .FF60_D1(w394), .ffxx(w395) );
	dmgcpu_WaveRAM waveram (.d[7](w103), .d[6](w104), .d[5](w105), .d[4](w106), .d[3](w107), .d[2](w108), .d[1](w109), .d[0](w110), .active(w376), .a[2](w377), .a[3](w378), .a[0](w379), .a[1](w380), .dout[0](w381), .dout[1](w382), .dout[2](w383), .dout[3](w384), .dout[4](w385), .dout[5](w386), .dout[6](w387), .dout[7](w388), .n_wr(w389), .bl_pch(w390), .n_rd(w391) );
	dmgcpu_and3 g1 (.a(1'b0), .b(w142) );
	dmgcpu_not g2 (.a(w370) );
endmodule // dmgcpu

// Module Definitions [It is possible to wrap here on your primitives]

module dmgcpu_IOBUF_B (  DRV_LOW, n_INPUT, n_ENA_PU, n_DRV_HIGH, PAD_IO);

	input wire DRV_LOW;
	output wire n_INPUT;
	input wire n_ENA_PU;
	input wire n_DRV_HIGH;
	inout wire PAD_IO;

endmodule // dmgcpu_IOBUF_B

module dmgcpu_IOBUF_C (  n_DRV_HIGH, n_ENA_PU, DRV_LOW, n_INPUT, PAD_IO);

	input wire n_DRV_HIGH;
	input wire n_ENA_PU;
	input wire DRV_LOW;
	output wire n_INPUT;
	inout wire PAD_IO;

endmodule // dmgcpu_IOBUF_C

module dmgcpu_IBUF_A (  n_INPUT, PAD_IN);

	output wire n_INPUT;
	input wire PAD_IN;

endmodule // dmgcpu_IBUF_A

module dmgcpu_IOBUF_A (  PAD_IO, n_DRV_HIGH, DRV_LOW, n_INPUT);

	inout wire PAD_IO;
	input wire n_DRV_HIGH;
	input wire DRV_LOW;
	output wire n_INPUT;

endmodule // dmgcpu_IOBUF_A

module dmgcpu_OBUF_A (  n_OUTPUT, PAD_OUT);

	input wire n_OUTPUT;
	output wire PAD_OUT;

endmodule // dmgcpu_OBUF_A

module dmgcpu_AOBUFFER (  VOUT, PAD_OUT);

	input wire VOUT;
	output wire PAD_OUT;

endmodule // dmgcpu_AOBUFFER

module dmgcpu_OBUF_B (  n_DRV_HIGH, DRV_LOW, PAD_OUT);

	input wire n_DRV_HIGH;
	input wire DRV_LOW;
	output wire PAD_OUT;

endmodule // dmgcpu_OBUF_B

module dmgcpu_IBUF_B (  PAD_IN, n_INPUT);

	input wire PAD_IN;
	output wire n_INPUT;

endmodule // dmgcpu_IBUF_B

module dmgcpu_OSC (  ENA, n_CLK, CK_IN, CK_OUT);

	input wire ENA;
	output wire n_CLK;
	input wire CK_IN;
	output wire CK_OUT;

endmodule // dmgcpu_OSC

module dmgcpu_AIBUFFER (  VIN, PAD_IN);

	output wire VIN;
	input wire PAD_IN;

endmodule // dmgcpu_AIBUFFER

module dmgcpu_PPU1 (  a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], n_ma[12], n_ma[10], n_ma[11], n_ma[8], n_ma[9], n_ma[6], n_ma[5], n_ma[7], n_ma[3], n_ma[2], n_ma[4], n_ma[1], n_ma[0], lcd_ld1, lcd_ld0, lcd_cpg, lcd_cp, lcd_st, lcd_cpl, lcd_fr, lcd_s, CONST0, n_dma_phi, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, ffxx, n_ppu_hard_reset, ff46, nma[9], fexx, nma[0], ff43, nma[4], nma[12], nma[6], nma[5], ff42, nma[11], nma[10], sprite_x_flip, nma[3], nma[2], sprite_x_match, bp_sel);

	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	output wire n_ma[12];
	output wire n_ma[10];
	output wire n_ma[11];
	output wire n_ma[8];
	output wire n_ma[9];
	output wire n_ma[6];
	output wire n_ma[5];
	output wire n_ma[7];
	output wire n_ma[3];
	output wire n_ma[2];
	output wire n_ma[4];
	output wire n_ma[1];
	output wire n_ma[0];
	output wire lcd_ld1;
	output wire lcd_ld0;
	output wire lcd_cpg;
	output wire lcd_cp;
	output wire lcd_st;
	output wire lcd_cpl;
	output wire lcd_fr;
	output wire lcd_s;
	input wire CONST0;
	input wire n_dma_phi;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire ppu_clk;
	input wire vram_to_oam;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	output wire ff46;
	inout wire nma[9];
	output wire fexx;
	inout wire nma[0];
	output wire ff43;
	inout wire nma[4];
	inout wire nma[12];
	inout wire nma[6];
	inout wire nma[5];
	output wire ff42;
	inout wire nma[11];
	inout wire nma[10];
	input wire sprite_x_flip;
	inout wire nma[3];
	inout wire nma[2];
	input wire sprite_x_match;
	output wire bp_sel;

endmodule // dmgcpu_PPU1

module dmgcpu_PPU2 (  cclk, clk6, n_reset2, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], n_oamb[0], n_oamb[1], n_oamb[2], n_oamb[3], n_oamb[4], n_oamb[5], n_oamb[6], n_oamb[7], oam_bl_pch, oa[1], oa[2], oa[3], oa[4], oa[5], oa[6], oa[7], n_oam_rd, n_oamb_wr, n_oama_wr, n_oama[0], n_oama[1], n_oama[2], n_oama[3], n_oama[4], n_oama[5], n_oama[6], n_oama[7], CONST0, n_dma_phi, dma_a[0], dma_a[4], dma_a[2], dma_a[6], dma_a[10], dma_a[1], dma_a[5], dma_a[11], dma_a[3], dma_a[7], dma_a[8], dma_a[12], dma_a[9], dma_run, soc_wr, soc_rd, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, n_ppu_hard_reset, nma[9], fexx, nma[0], ff43, nma[4], nma[12], nma[6], nma[5], ff42, nma[11], nma[10], sprite_x_flip, nma[3], nma[2], sprite_x_match, bp_sel);

	input wire cclk;
	input wire clk6;
	input wire n_reset2;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	inout wire n_oamb[0];
	inout wire n_oamb[1];
	inout wire n_oamb[2];
	inout wire n_oamb[3];
	inout wire n_oamb[4];
	inout wire n_oamb[5];
	inout wire n_oamb[6];
	inout wire n_oamb[7];
	output wire oam_bl_pch;
	output wire oa[1];
	output wire oa[2];
	output wire oa[3];
	output wire oa[4];
	output wire oa[5];
	output wire oa[6];
	output wire oa[7];
	output wire n_oam_rd;
	output wire n_oamb_wr;
	output wire n_oama_wr;
	inout wire n_oama[0];
	inout wire n_oama[1];
	inout wire n_oama[2];
	inout wire n_oama[3];
	inout wire n_oama[4];
	inout wire n_oama[5];
	inout wire n_oama[6];
	inout wire n_oama[7];
	input wire CONST0;
	input wire n_dma_phi;
	input wire dma_a[0];
	input wire dma_a[4];
	input wire dma_a[2];
	input wire dma_a[6];
	input wire dma_a[10];
	input wire dma_a[1];
	input wire dma_a[5];
	input wire dma_a[11];
	input wire dma_a[3];
	input wire dma_a[7];
	input wire dma_a[8];
	input wire dma_a[12];
	input wire dma_a[9];
	input wire dma_run;
	input wire soc_wr;
	input wire soc_rd;
	output wire ppu_rd;
	output wire ppu_wr;
	output wire ppu_clk;
	input wire vram_to_oam;
	output wire n_ppu_hard_reset;
	inout wire nma[9];
	input wire fexx;
	inout wire nma[0];
	input wire ff43;
	inout wire nma[4];
	inout wire nma[12];
	inout wire nma[6];
	inout wire nma[5];
	input wire ff42;
	inout wire nma[11];
	inout wire nma[10];
	output wire sprite_x_flip;
	inout wire nma[3];
	inout wire nma[2];
	output wire sprite_x_match;
	input wire bp_sel;

endmodule // dmgcpu_PPU2

module dmgcpu_OAM (  n_oamb[0], n_oamb[1], n_oamb[2], n_oamb[3], n_oamb[4], n_oamb[5], n_oamb[6], n_oamb[7], oam_bl_pch, oa[1], oa[2], oa[3], oa[4], oa[5], oa[6], oa[7], n_oam_rd, n_oamb_wr, n_oama_wr, n_oama[0], n_oama[1], n_oama[2], n_oama[3], n_oama[4], n_oama[5], n_oama[6], n_oama[7]);

	inout wire n_oamb[0];
	inout wire n_oamb[1];
	inout wire n_oamb[2];
	inout wire n_oamb[3];
	inout wire n_oamb[4];
	inout wire n_oamb[5];
	inout wire n_oamb[6];
	inout wire n_oamb[7];
	input wire oam_bl_pch;
	input wire oa[1];
	input wire oa[2];
	input wire oa[3];
	input wire oa[4];
	input wire oa[5];
	input wire oa[6];
	input wire oa[7];
	input wire n_oam_rd;
	input wire n_oamb_wr;
	input wire n_oama_wr;
	inout wire n_oama[0];
	inout wire n_oama[1];
	inout wire n_oama[2];
	inout wire n_oama[3];
	inout wire n_oama[4];
	inout wire n_oama[5];
	inout wire n_oama[6];
	inout wire n_oama[7];

endmodule // dmgcpu_OAM

module dmgcpu_HRAM (  clk7, a[0], a[1], d[7], d[6], d[5], d[4, d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], soc_wr, soc_rd, ffxx);

	input wire clk7;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4;
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire soc_wr;
	input wire soc_rd;
	input wire ffxx;

endmodule // dmgcpu_HRAM

module dmgcpu_DAC (  vin_analog, so2_analog, so1_analog);

	input wire vin_analog;
	output wire so2_analog;
	output wire so1_analog;

endmodule // dmgcpu_DAC

module dmgcpu_BootROM (  a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15]);

	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	input wire a[15];

endmodule // dmgcpu_BootROM

module dmgcpu_Ser (  n_reset2, d[5], d[6], d[7], d[4], d[3], d[2], d[1], d[0], n_sin, sck_dir, n_sck, int_serial, sc_read, sb_read, sc_write, n_sb_write, lfo_16384Hz, ser_out, serial_tick);

	input wire n_reset2;
	inout wire d[5];
	inout wire d[6];
	inout wire d[7];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire n_sin;
	output wire sck_dir;
	input wire n_sck;
	output wire int_serial;
	input wire sc_read;
	input wire sb_read;
	input wire sc_write;
	input wire n_sb_write;
	input wire lfo_16384Hz;
	output wire ser_out;
	output wire serial_tick;

endmodule // dmgcpu_Ser

module dmgcpu_ClkGen (  n_clk_in, reset, cclk, clk1, clk2, clk3, clk4, osc_stable, clk_ena, osc_ena, clk5, clk6, clk7, clk8, clk9, n_reset2, sync_reset, cpu_mreq, ext_cs_en, cpu_wr_sync, cpu_wr, test_1, n_test_reset);

	input wire n_clk_in;
	input wire reset;
	output wire cclk;
	output wire clk1;
	output wire clk2;
	output wire clk3;
	output wire clk4;
	input wire osc_stable;
	input wire clk_ena;
	input wire osc_ena;
	output wire clk5;
	output wire clk6;
	output wire clk7;
	output wire clk8;
	output wire clk9;
	output wire n_reset2;
	output wire sync_reset;
	input wire cpu_mreq;
	output wire ext_cs_en;
	output wire cpu_wr_sync;
	input wire cpu_wr;
	input wire test_1;
	input wire n_test_reset;

endmodule // dmgcpu_ClkGen

module dmgcpu_MMIO (  reset, clk2, clk4, osc_stable, clk_ena, osc_ena, clk6, clk9, n_reset2, cpu_wr_sync, cpu_m1, n_cpu_m1, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], cpu_irq_trig[4], cpu_irq_ack[4], cpu_irq_trig[3], cpu_irq_ack[3], cpu_irq_trig[2], cpu_irq_ack[2], cpu_irq_trig[1], cpu_irq_ack[1], cpu_irq_trig[0], cpu_irq_ack[0], cpu_rd, cpu_wr, n_DRV_HIGH_a[14], n_INPUT_a[14], DRV_LOW_a[14], n_DRV_HIGH_a[13], n_INPUT_a[13], DRV_LOW_a[13], n_DRV_HIGH_a[12], n_INPUT_a[12], DRV_LOW_a[12], n_DRV_HIGH_a[11], n_INPUT_a[11], DRV_LOW_a[11], n_DRV_HIGH_a[10], n_INPUT_a[10], DRV_LOW_a[10], n_DRV_HIGH_a[9], n_INPUT_a[9], DRV_LOW_a[9], n_DRV_HIGH_a[8], n_INPUT_a[8], DRV_LOW_a[8], n_DRV_HIGH_nrd, n_INPUT_nrd, DRV_LOW_nrd, n_DRV_HIGH_nwr, n_INPUT_nwr, DRV_LOW_nwr, n_t1_frompad, n_t2_frompad, CONST0, n_ena_pu_db, n_dma_phi, dma_a[0], dma_a[4], dma_a[2], dma_a[6], dma_a[10], dma_a[1], dma_a[5], dma_a[11], dma_a[3], dma_a[7], dma_a[8], dma_a[12], dma_a[9], dma_run, soc_wr, soc_rd, lfo_512Hz, ppu_rd, ppu_wr, int_serial, sc_read, sb_read, sc_write, n_sb_write, lfo_16384Hz, ppu_clk, vram_to_oam, dma_a[15], non_vram_mreq, test_1, test_2, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, n_test_reset, n_ext_addr_en, addr_latch, int_jp, FF60_D1, ffxx, n_ppu_hard_reset, ff46);

	input wire reset;
	input wire clk2;
	input wire clk4;
	output wire osc_stable;
	input wire clk_ena;
	input wire osc_ena;
	input wire clk6;
	input wire clk9;
	input wire n_reset2;
	input wire cpu_wr_sync;
	input wire cpu_m1;
	output wire n_cpu_m1;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	output wire cpu_irq_trig[4];
	input wire cpu_irq_ack[4];
	output wire cpu_irq_trig[3];
	input wire cpu_irq_ack[3];
	output wire cpu_irq_trig[2];
	input wire cpu_irq_ack[2];
	output wire cpu_irq_trig[1];
	input wire cpu_irq_ack[1];
	output wire cpu_irq_trig[0];
	input wire cpu_irq_ack[0];
	input wire cpu_rd;
	input wire cpu_wr;
	output wire n_DRV_HIGH_a[14];
	input wire n_INPUT_a[14];
	output wire DRV_LOW_a[14];
	output wire n_DRV_HIGH_a[13];
	input wire n_INPUT_a[13];
	output wire DRV_LOW_a[13];
	output wire n_DRV_HIGH_a[12];
	input wire n_INPUT_a[12];
	output wire DRV_LOW_a[12];
	output wire n_DRV_HIGH_a[11];
	input wire n_INPUT_a[11];
	output wire DRV_LOW_a[11];
	output wire n_DRV_HIGH_a[10];
	input wire n_INPUT_a[10];
	output wire DRV_LOW_a[10];
	output wire n_DRV_HIGH_a[9];
	input wire n_INPUT_a[9];
	output wire DRV_LOW_a[9];
	output wire n_DRV_HIGH_a[8];
	input wire n_INPUT_a[8];
	output wire DRV_LOW_a[8];
	output wire n_DRV_HIGH_nrd;
	input wire n_INPUT_nrd;
	output wire DRV_LOW_nrd;
	output wire n_DRV_HIGH_nwr;
	input wire n_INPUT_nwr;
	output wire DRV_LOW_nwr;
	input wire n_t1_frompad;
	input wire n_t2_frompad;
	input wire CONST0;
	output wire n_ena_pu_db;
	output wire n_dma_phi;
	output wire dma_a[0];
	output wire dma_a[4];
	output wire dma_a[2];
	output wire dma_a[6];
	output wire dma_a[10];
	output wire dma_a[1];
	output wire dma_a[5];
	output wire dma_a[11];
	output wire dma_a[3];
	output wire dma_a[7];
	output wire dma_a[8];
	output wire dma_a[12];
	output wire dma_a[9];
	output wire dma_run;
	output wire soc_wr;
	output wire soc_rd;
	output wire lfo_512Hz;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire int_serial;
	output wire sc_read;
	output wire sb_read;
	output wire sc_write;
	output wire n_sb_write;
	output wire lfo_16384Hz;
	input wire ppu_clk;
	output wire vram_to_oam;
	output wire dma_a[15];
	input wire non_vram_mreq;
	output wire test_1;
	output wire test_2;
	output wire n_extdb_to_intdb;
	output wire n_dblatch_to_intdb;
	output wire n_intdb_to_extdb;
	output wire n_test_reset;
	output wire n_ext_addr_en;
	output wire addr_latch;
	input wire int_jp;
	input wire FF60_D1;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ff46;

endmodule // dmgcpu_MMIO

module dmgcpu_SM83Core (  RESET, CLK1, CLK2, CLK3, CLK4, OSC_STABLE, CLK_ENA, OSC_ENA, CLK5, CLK6, CLK7, CLK8, CLK9, SYNC_RESET, CPU_MREQ, NMI, M1, A[0], A[1], D[7], D[6], D[5], D[4], D[3], D[2], D[1], D[0], A[2], A[3], A[4], A[5], A[6], A[7], A[8], A[9], A[10], A[11], A[12], A[13], A[14], A[15], CPU_IRQ_TRIG[7], CPU_IRQ_ACK[7], CPU_IRQ_TRIG[6], CPU_IRQ_ACK[6], CPU_IRQ_TRIG[5], CPU_IRQ_ACK[5], CPU_IRQ_TRIG[4], CPU_IRQ_ACK[4], CPU_IRQ_TRIG[3], CPU_IRQ_ACK[3], CPU_IRQ_TRIG[2], CPU_IRQ_ACK[2], CPU_IRQ_TRIG[1], CPU_IRQ_ACK[1], CPU_IRQ_TRIG[0], CPU_IRQ_ACK[0], WAKE, RD, WR, MMIO_REQ, IPL_REQ, BUS_DISABLE, IPL_DISABLE);

	input wire RESET;
	input wire CLK1;
	input wire CLK2;
	input wire CLK3;
	input wire CLK4;
	input wire OSC_STABLE;
	output wire CLK_ENA;
	output wire OSC_ENA;
	input wire CLK5;
	input wire CLK6;
	input wire CLK7;
	input wire CLK8;
	input wire CLK9;
	input wire SYNC_RESET;
	output wire CPU_MREQ;
	input wire NMI;
	output wire M1;
	output wire A[0];
	output wire A[1];
	inout wire D[7];
	inout wire D[6];
	inout wire D[5];
	inout wire D[4];
	inout wire D[3];
	inout wire D[2];
	inout wire D[1];
	inout wire D[0];
	output wire A[2];
	output wire A[3];
	output wire A[4];
	output wire A[5];
	output wire A[6];
	output wire A[7];
	output wire A[8];
	output wire A[9];
	output wire A[10];
	output wire A[11];
	output wire A[12];
	output wire A[13];
	output wire A[14];
	output wire A[15];
	input wire CPU_IRQ_TRIG[7];
	output wire CPU_IRQ_ACK[7];
	input wire CPU_IRQ_TRIG[6];
	output wire CPU_IRQ_ACK[6];
	input wire CPU_IRQ_TRIG[5];
	output wire CPU_IRQ_ACK[5];
	input wire CPU_IRQ_TRIG[4];
	output wire CPU_IRQ_ACK[4];
	input wire CPU_IRQ_TRIG[3];
	output wire CPU_IRQ_ACK[3];
	input wire CPU_IRQ_TRIG[2];
	output wire CPU_IRQ_ACK[2];
	input wire CPU_IRQ_TRIG[1];
	output wire CPU_IRQ_ACK[1];
	input wire CPU_IRQ_TRIG[0];
	output wire CPU_IRQ_ACK[0];
	input wire WAKE;
	output wire RD;
	output wire WR;
	input wire MMIO_REQ;
	input wire IPL_REQ;
	input wire BUS_DISABLE;
	input wire IPL_DISABLE;

endmodule // dmgcpu_SM83Core

module dmgcpu_Arbiter (  clk2, n_reset2, cpu_mreq, ext_cs_en, cpu_wr_sync, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], cpu_wr, mmio_sel, boot_sel, n_DRV_HIGH_a[15], n_INPUT_a[15], DRV_LOW_a[15], n_cs_topad, CONST0, n_DRV_HIGH_nmwr, n_mwr, DRV_LOW_nmwr, n_DRV_HIGH_nmrd, n_mrd, DRV_LOW_nmrd, n_DRV_HIGH_nmcs, n_mcs, DRV_LOW_nmcs, n_DRV_HIGH_md[7], n_md_frompad[7], DRV_LOW_md[7], n_md_ena_pu, n_DRV_HIGH_md[6], n_md_frompad[6], DRV_LOW_md[6], n_DRV_HIGH_md[5], n_md_frompad[5], DRV_LOW_md[5], n_DRV_HIGH_md[4], n_md_frompad[4], DRV_LOW_md[4], n_DRV_HIGH_md[3], n_md_frompad[3], DRV_LOW_md[3], n_DRV_HIGH_md[2], n_md_frompad[2], DRV_LOW_md[2], n_DRV_HIGH_md[1], n_md_frompad[1], DRV_LOW_md[1], n_DRV_HIGH_md[0], DRV_LOW_md[0], n_md_frompad[0], n_DRV_HIGH_d[7], n_db_frompad[7], DRV_LOW_d[7], n_ena_pu_db, n_DRV_HIGH_d[6], n_db_frompad[6], DRV_LOW_d[6], n_DRV_HIGH_d[5], n_db_frompad[5], DRV_LOW_d[5], n_DRV_HIGH_d[4], n_db_frompad[4], DRV_LOW_d[4], n_DRV_HIGH_d[3], n_db_frompad[3], DRV_LOW_d[3], n_DRV_HIGH_d[2], n_db_frompad[2], DRV_LOW_d[2], n_DRV_HIGH_d[1], n_db_frompad[1], DRV_LOW_d[1], n_DRV_HIGH_d[0], n_db_frompad[0], DRV_LOW_a[0], soc_wr, soc_rd, vram_to_oam, dma_a[15], non_vram_mreq, test_1, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, ffxx, n_ppu_hard_reset);

	input wire clk2;
	input wire n_reset2;
	input wire cpu_mreq;
	input wire ext_cs_en;
	input wire cpu_wr_sync;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	input wire a[15];
	input wire cpu_wr;
	output wire mmio_sel;
	output wire boot_sel;
	output wire n_DRV_HIGH_a[15];
	input wire n_INPUT_a[15];
	output wire DRV_LOW_a[15];
	output wire n_cs_topad;
	output wire CONST0;
	output wire n_DRV_HIGH_nmwr;
	input wire n_mwr;
	output wire DRV_LOW_nmwr;
	output wire n_DRV_HIGH_nmrd;
	input wire n_mrd;
	output wire DRV_LOW_nmrd;
	output wire n_DRV_HIGH_nmcs;
	input wire n_mcs;
	output wire DRV_LOW_nmcs;
	output wire n_DRV_HIGH_md[7];
	input wire n_md_frompad[7];
	output wire DRV_LOW_md[7];
	output wire n_md_ena_pu;
	output wire n_DRV_HIGH_md[6];
	input wire n_md_frompad[6];
	output wire DRV_LOW_md[6];
	output wire n_DRV_HIGH_md[5];
	input wire n_md_frompad[5];
	output wire DRV_LOW_md[5];
	output wire n_DRV_HIGH_md[4];
	input wire n_md_frompad[4];
	output wire DRV_LOW_md[4];
	output wire n_DRV_HIGH_md[3];
	input wire n_md_frompad[3];
	output wire DRV_LOW_md[3];
	output wire n_DRV_HIGH_md[2];
	input wire n_md_frompad[2];
	output wire DRV_LOW_md[2];
	output wire n_DRV_HIGH_md[1];
	input wire n_md_frompad[1];
	output wire DRV_LOW_md[1];
	output wire n_DRV_HIGH_md[0];
	output wire DRV_LOW_md[0];
	input wire n_md_frompad[0];
	output wire n_DRV_HIGH_d[7];
	input wire n_db_frompad[7];
	output wire DRV_LOW_d[7];
	input wire n_ena_pu_db;
	output wire n_DRV_HIGH_d[6];
	input wire n_db_frompad[6];
	output wire DRV_LOW_d[6];
	output wire n_DRV_HIGH_d[5];
	input wire n_db_frompad[5];
	output wire DRV_LOW_d[5];
	output wire n_DRV_HIGH_d[4];
	input wire n_db_frompad[4];
	output wire DRV_LOW_d[4];
	output wire n_DRV_HIGH_d[3];
	input wire n_db_frompad[3];
	output wire DRV_LOW_d[3];
	output wire n_DRV_HIGH_d[2];
	input wire n_db_frompad[2];
	output wire DRV_LOW_d[2];
	output wire n_DRV_HIGH_d[1];
	input wire n_db_frompad[1];
	output wire DRV_LOW_d[1];
	output wire n_DRV_HIGH_d[0];
	input wire n_db_frompad[0];
	output wire DRV_LOW_a[0];
	input wire soc_wr;
	input wire soc_rd;
	input wire vram_to_oam;
	input wire dma_a[15];
	output wire non_vram_mreq;
	input wire test_1;
	input wire n_extdb_to_intdb;
	input wire n_dblatch_to_intdb;
	input wire n_intdb_to_extdb;
	output wire ffxx;
	input wire n_ppu_hard_reset;

endmodule // dmgcpu_Arbiter

module dmgcpu_APU (  cclk, clk2, clk4, clk6, clk7, clk9, n_reset2, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], cpu_wakeup, n_DRV_HIGH_a[7], n_INPUT_a[7], DRV_LOW_a[7], n_DRV_HIGH_a[6], n_INPUT_a[6], DRV_LOW_a[6], n_DRV_HIGH_a[5], n_INPUT_a[5], DRV_LOW_a[5], n_DRV_HIGH_a[4], n_INPUT_a[4], DRV_LOW_a[4], n_DRV_HIGH_a[3], n_INPUT_a[3], DRV_LOW_a[3], n_DRV_HIGH_a[2], n_INPUT_a[2], DRV_LOW_a[2], n_DRV_HIGH_a[1], n_INPUT_a[1], DRV_LOW_a[1], n_DRV_HIGH_a[0], n_INPUT_a[0], DRV_LOW_a[0], n_sout_topad, n_DRV_HIGH_sin, n_ENA_PU_sin, DRV_LOW_sin, n_DRV_HIGH_sck, sck_dir, DRV_LOW_sck, n_DRV_HIGH_p10, CONST0, n_p10, DRV_LOW_p10, n_DRV_HIGH_p11, n_p11, DRV_LOW_p11, n_DRV_HIGH_p12, n_p12, DRV_LOW_p12, n_DRV_HIGH_p13, n_p13, DRV_LOW_p13, n_DRV_HIGH_p14, DRV_LOW_p14, n_DRV_HIGH_p15, DRV_LOW_p15, dma_a[0], dma_a[4], dma_a[2], dma_a[6], dma_a[1], dma_a[5], dma_a[3], dma_a[7], soc_wr, soc_rd, lfo_512Hz, ser_out, serial_tick, test_1, test_2, n_ext_addr_en, ch3_active, wave_a[2], wave_a[3], wave_a[0], wave_a[1], wave_rd[0], wave_rd[1], wave_rd[2], wave_rd[3], wave_rd[4], wave_rd[5], wave_rd[6], wave_rd[7], n_wave_wr, wave_bl_pch, n_wave_rd, addr_latch, int_jp, FF60_D1, ffxx);

	input wire cclk;
	input wire clk2;
	input wire clk4;
	input wire clk6;
	input wire clk7;
	input wire clk9;
	input wire n_reset2;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	output wire cpu_wakeup;
	output wire n_DRV_HIGH_a[7];
	input wire n_INPUT_a[7];
	output wire DRV_LOW_a[7];
	output wire n_DRV_HIGH_a[6];
	input wire n_INPUT_a[6];
	output wire DRV_LOW_a[6];
	output wire n_DRV_HIGH_a[5];
	input wire n_INPUT_a[5];
	output wire DRV_LOW_a[5];
	output wire n_DRV_HIGH_a[4];
	input wire n_INPUT_a[4];
	output wire DRV_LOW_a[4];
	output wire n_DRV_HIGH_a[3];
	input wire n_INPUT_a[3];
	output wire DRV_LOW_a[3];
	output wire n_DRV_HIGH_a[2];
	input wire n_INPUT_a[2];
	output wire DRV_LOW_a[2];
	output wire n_DRV_HIGH_a[1];
	input wire n_INPUT_a[1];
	output wire DRV_LOW_a[1];
	output wire n_DRV_HIGH_a[0];
	input wire n_INPUT_a[0];
	output wire DRV_LOW_a[0];
	output wire n_sout_topad;
	output wire n_DRV_HIGH_sin;
	output wire n_ENA_PU_sin;
	output wire DRV_LOW_sin;
	output wire n_DRV_HIGH_sck;
	input wire sck_dir;
	output wire DRV_LOW_sck;
	output wire n_DRV_HIGH_p10;
	input wire CONST0;
	input wire n_p10;
	output wire DRV_LOW_p10;
	output wire n_DRV_HIGH_p11;
	input wire n_p11;
	output wire DRV_LOW_p11;
	output wire n_DRV_HIGH_p12;
	input wire n_p12;
	output wire DRV_LOW_p12;
	output wire n_DRV_HIGH_p13;
	input wire n_p13;
	output wire DRV_LOW_p13;
	output wire n_DRV_HIGH_p14;
	output wire DRV_LOW_p14;
	output wire n_DRV_HIGH_p15;
	output wire DRV_LOW_p15;
	input wire dma_a[0];
	input wire dma_a[4];
	input wire dma_a[2];
	input wire dma_a[6];
	input wire dma_a[1];
	input wire dma_a[5];
	input wire dma_a[3];
	input wire dma_a[7];
	input wire soc_wr;
	input wire soc_rd;
	input wire lfo_512Hz;
	input wire ser_out;
	input wire serial_tick;
	input wire test_1;
	input wire test_2;
	input wire n_ext_addr_en;
	output wire ch3_active;
	output wire wave_a[2];
	output wire wave_a[3];
	output wire wave_a[0];
	output wire wave_a[1];
	input wire wave_rd[0];
	input wire wave_rd[1];
	input wire wave_rd[2];
	input wire wave_rd[3];
	input wire wave_rd[4];
	input wire wave_rd[5];
	input wire wave_rd[6];
	input wire wave_rd[7];
	output wire n_wave_wr;
	output wire wave_bl_pch;
	output wire n_wave_rd;
	input wire addr_latch;
	output wire int_jp;
	output wire FF60_D1;
	input wire ffxx;

endmodule // dmgcpu_APU

module dmgcpu_WaveRAM (  d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], active, a[2], a[3], a[0], a[1], dout[0], dout[1], dout[2], dout[3], dout[4], dout[5], dout[6], dout[7], n_wr, bl_pch, n_rd);

	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire active;
	input wire a[2];
	input wire a[3];
	input wire a[0];
	input wire a[1];
	output wire dout[0];
	output wire dout[1];
	output wire dout[2];
	output wire dout[3];
	output wire dout[4];
	output wire dout[5];
	output wire dout[6];
	output wire dout[7];
	input wire n_wr;
	input wire bl_pch;
	input wire n_rd;

endmodule // dmgcpu_WaveRAM

module dmgcpu_and3 (  a, b, c, x);

	input wire a;
	input wire b;
	input wire c;
	output wire x;

endmodule // dmgcpu_and3

module dmgcpu_not (  a, x);

	input wire a;
	output wire x;

endmodule // dmgcpu_not



// ERROR: floating wire w125
// ERROR: floating wire w126
// ERROR: floating wire w127
// ERROR: floating wire w143
// WARNING: wire not driving anything w286
// WARNING: wire not driving anything w336
// WARNING: Cell dmgcpu_IOBUF_B:pad_d0 port DRV_LOW not connected.
// WARNING: Cell dmgcpu_IOBUF_A:pad_nmcs port DRV_LOW not connected.
// WARNING: Cell dmgcpu_OBUF_A:pad_m1 port PAD_OUT not connected.
// WARNING: Cell dmgcpu_IBUF_B:pad_nnmi port PAD_IN not connected.
// WARNING: Cell dmgcpu_SM83Core:core port CPU_IRQ_ACK[7] not connected.
// WARNING: Cell dmgcpu_SM83Core:core port CPU_IRQ_ACK[6] not connected.
// WARNING: Cell dmgcpu_SM83Core:core port CPU_IRQ_ACK[5] not connected.
// WARNING: Cell dmgcpu_and3:g1 port c not connected.
// WARNING: Cell dmgcpu_and3:g1 port x not connected.
// WARNING: Cell dmgcpu_not:g2 port x not connected.
