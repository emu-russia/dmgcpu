
module Decoder1 (CLK, a, d);

	input CLK;
	input [25:0] a;
	output [106:0] d;

endmodule // Decoder1
