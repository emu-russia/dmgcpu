module BootROM (  a, d, from_g1_YULA);

	input wire [15:0] a;
	inout wire [7:0] d;
	input wire from_g1_YULA;

endmodule // BootROM