module MMIO (  reset, clk2, clk4, osc_stable, clk_ena, osc_ena, clk6, clk9, n_reset2, cpu_wr_sync, cpu_m1, n_cpu_m1, 
	a, d, 
	cpu_irq_trig, cpu_irq_ack, cpu_rd, cpu_wr, 
	n_DRV_HIGH_a, n_INPUT_a, DRV_LOW_a, 
	n_DRV_HIGH_nrd, n_INPUT_nrd, DRV_LOW_nrd, n_DRV_HIGH_nwr, n_INPUT_nwr, DRV_LOW_nwr, n_t1_frompad, n_t2_frompad, CONST0, n_ena_pu_db, n_dma_phi, 
	dma_a, dma_a_15, dma_run, soc_wr, soc_rd, lfo_512Hz, ppu_rd, ppu_wr, int_serial, sc_read, sb_read, sc_write, n_sb_write, lfo_16384Hz, ppu_clk, vram_to_oam, non_vram_mreq, 
	test_1, test_2, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, n_test_reset, n_ext_addr_en, addr_latch, int_jp, FF60_D1, ffxx, n_ppu_hard_reset, ff46, dma_addr_ext, cpu_vram_oam_rd, oam_dma_wr, ppu_int_stat, ppu_int_vbl, clk6_delay);

	input wire reset;
	input wire clk2;
	input wire clk4;
	output wire osc_stable;
	input wire clk_ena;
	input wire osc_ena;
	input wire clk6;
	input wire clk9;
	input wire n_reset2;
	input wire cpu_wr_sync;
	input wire cpu_m1;
	output wire n_cpu_m1;
	inout wire [14:0] a; 			// a[15] is not used    ⚠️ bidir
	inout wire [7:0] d;
	output wire [4:0] cpu_irq_trig;
	input wire [4:0] cpu_irq_ack;
	input wire cpu_rd;
	input wire cpu_wr;
	output wire [14:8] n_DRV_HIGH_a;
	input wire [14:8] n_INPUT_a;
	output wire [14:8] DRV_LOW_a;
	output wire n_DRV_HIGH_nrd;
	input wire n_INPUT_nrd;
	output wire DRV_LOW_nrd;
	output wire n_DRV_HIGH_nwr;
	input wire n_INPUT_nwr;
	output wire DRV_LOW_nwr;
	input wire n_t1_frompad;
	input wire n_t2_frompad;
	inout wire CONST0;
	output wire n_ena_pu_db;
	output wire n_dma_phi;
	output wire [12:0] dma_a;
	output wire dma_a_15;
	output wire dma_run;
	output wire soc_wr;
	output wire soc_rd;
	output wire lfo_512Hz;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire int_serial;
	output wire sc_read;
	output wire sb_read;
	output wire sc_write;
	output wire n_sb_write;
	output wire lfo_16384Hz;
	input wire ppu_clk;
	output wire vram_to_oam;
	input wire non_vram_mreq;
	output wire test_1;
	output wire test_2;
	output wire n_extdb_to_intdb;
	output wire n_dblatch_to_intdb;
	output wire n_intdb_to_extdb;
	output wire n_test_reset;
	output wire n_ext_addr_en;
	output wire addr_latch;
	input wire int_jp;
	input wire FF60_D1;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ff46;
	output wire dma_addr_ext;
	output wire cpu_vram_oam_rd;
	output wire oam_dma_wr;
	input wire ppu_int_stat;
	input wire ppu_int_vbl;
	input wire clk6_delay;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;

	assign DRV_LOW_a[13] = w1;
	assign n_DRV_HIGH_a[13] = w7;
	assign w6 = n_INPUT_a[13];
	assign n_DRV_HIGH_a[12] = w51;
	assign DRV_LOW_a[12] = w291;
	assign n_DRV_HIGH_a[11] = w290;
	assign w235 = n_INPUT_a[8];
	assign n_DRV_HIGH_a[9] = w236;
	assign DRV_LOW_a[9] = w270;
	assign n_DRV_HIGH_a[8] = w293;
	assign DRV_LOW_a[8] = w294;
	assign w10 = n_INPUT_a[11];
	assign DRV_LOW_a[11] = w292;
	assign w269 = n_INPUT_a[9];
	assign w264 = clk_ena;
	assign w265 = n_INPUT_a[14];
	assign n_DRV_HIGH_a[14] = w267;
	assign DRV_LOW_a[14] = w268;
	assign osc_stable = w364;
	assign DRV_LOW_a[10] = w289;
	assign n_DRV_HIGH_a[10] = w34;
	assign w213 = n_INPUT_a[10];
	assign w358 = int_serial;
	assign test_2 = w215;
	assign n_test_reset = w54;
	assign lfo_16384Hz = w53;
	assign sc_write = w317;
	assign w160 = n_INPUT_nrd;
	assign sc_read = w146;
	assign n_DRV_HIGH_nrd = w35;
	assign sb_read = w145;
	assign w74 = clk9;
	assign n_ext_addr_en = w8;
	assign DRV_LOW_nwr = w216;
	assign w217 = n_INPUT_nwr;
	assign DRV_LOW_nrd = w41;
	assign n_DRV_HIGH_nwr = w40;
	assign n_sb_write = w359;
	assign w39 = n_t1_frompad;
	assign w52 = n_t2_frompad;
	assign w63 = n_reset2;
	assign addr_latch = w130;
	assign w86 = int_jp;
	assign w87 = FF60_D1;
	assign test_1 = w36;
	assign dma_addr_ext = w89;
	assign w312 = clk4;
	assign lfo_512Hz = w113;
	assign a[0] = w112;
	assign soc_wr = w110;
	assign a[1] = w108;
	assign a[3] = w249;
	assign a[5] = w107;
	assign a[6] = w250;
	assign a[2] = w306;
	assign a[7] = w251;
	assign a[4] = w103;
	assign d[1] = w68;
	assign d[2] = w71;
	assign d[0] = w31;
	assign d[6] = w118;
	assign d[5] = w19;
	assign d[3] = w23;
	assign d[4] = w95;
	assign d[7] = w155;
	assign soc_rd = w45;
	assign CONST0 = w20;
	assign dma_a[5] = w281;
	assign dma_a[1] = w173;
	assign dma_a[6] = w172;
	assign dma_a[3] = w343;
	assign n_cpu_m1 = w287;
	assign dma_a[2] = w247;
	assign w148 = ffxx;
	assign dma_a[0] = w174;
	assign dma_a[4] = w175;
	assign oam_dma_wr = w344;
	assign dma_a[10] = w282;
	assign dma_a[7] = w179;
	assign w180 = ppu_clk;
	assign w206 = clk6;
	assign dma_a[11] = w207;
	assign w241 = ppu_wr;
	assign w184 = clk6_delay;
	assign dma_a[12] = w158;
	assign dma_run = w185;
	assign w240 = ff46;
	assign dma_a[8] = w239;
	assign n_dma_phi = w323;
	assign w188 = n_ppu_hard_reset;
	assign dma_a[9] = w276;
	assign w286 = cpu_m1;
	assign cpu_vram_oam_rd = w182;
	assign cpu_irq_trig[4] = w131;
	assign w259 = ppu_int_stat;
	assign w132 = cpu_irq_ack[4];
	assign a[10] = w320;
	assign w260 = clk2;
	assign w168 = cpu_irq_ack[3];
	assign vram_to_oam = w169;
	assign w65 = ppu_int_vbl;
	assign w257 = cpu_irq_ack[2];
	assign cpu_irq_trig[1] = w152;
	assign cpu_irq_trig[2] = w153;
	assign cpu_irq_trig[3] = w162;
	assign w163 = cpu_irq_ack[1];
	assign cpu_irq_trig[0] = w164;
	assign w324 = cpu_irq_ack[0];
	assign w263 = non_vram_mreq;
	assign dma_a_15 = w192;
	assign w202 = osc_ena;
	assign a[13] = w4;
	assign w201 = cpu_wr;
	assign n_extdb_to_intdb = w302;
	assign n_dblatch_to_intdb = w262;
	assign w55 = reset;
	assign n_intdb_to_extdb = w261;
	assign w203 = cpu_wr_sync;
	assign a[14] = w28;
	assign n_ena_pu_db = w299;
	assign a[11] = w48;
	assign w47 = cpu_rd;
	assign a[8] = w272;
	assign a[9] = w229;
	assign a[12] = w49;
	assign w295 = n_INPUT_a[12];

	// Instances

	dmg_not g1 (.a(w6), .x(w5) );
	dmg_not g2 (.a(w295), .x(w50) );
	dmg_not g3 (.a(w275), .x(w274) );
	dmg_not g4 (.a(w200), .x(w199) );
	dmg_not g5 (.a(w263), .x(w325) );
	dmg_not g6 (.a(w324), .x(w193) );
	dmg_not g7 (.a(w261), .x(w299) );
	dmg_not g8 (.a(w192), .x(w191) );
	dmg_not g9 (.a(w163), .x(w66) );
	dmg_not g10 (.a(w170), .x(w169) );
	dmg_not g11 (.a(w257), .x(w256) );
	dmg_not g12 (.a(w168), .x(w167) );
	dmg_not g13 (.a(w132), .x(w70) );
	dmg_not g14 (.a(w285), .x(w177) );
	dmg_not g15 (.a(w190), .x(w284) );
	dmg_not g16 (.a(w283), .x(w89) );
	dmg_not g17 (.a(w242), .x(w243) );
	dmg_not g18 (.a(w286), .x(w287) );
	dmg_not g19 (.a(w310), .x(w309) );
	dmg_not g20 (.a(w341), .x(w342) );
	dmg_not g21 (.a(w269), .x(w11) );
	dmg_not g22 (.a(w116), .x(w117) );
	dmg_not g23 (.a(w32), .x(w69) );
	dmg_not g24 (.a(w45), .x(w44) );
	dmg_not g25 (.a(w137), .x(w138) );
	dmg_not g26 (.a(w36), .x(w8) );
	dmg_not g27 (.a(w141), .x(w140) );
	dmg_not g28 (.a(w39), .x(w38) );
	dmg_not g29 (.a(w52), .x(w161) );
	dmg_not g30 (.a(w219), .x(w53) );
	dmg_not g31 (.a(w202), .x(w56) );
	dmg_not g32 (.a(w143), .x(w144) );
	dmg_not g33 (.a(w79), .x(w78) );
	dmg_not g34 (.a(w81), .x(w82) );
	dmg_not g35 (.a(w314), .x(w313) );
	dmg_not g36 (.a(w114), .x(w113) );
	dmg_not g37 (.a(w105), .x(w106) );
	dmg_not g38 (.a(w306), .x(w305) );
	dmg_not g39 (.a(w315), .x(w345) );
	dmg_not g40 (.a(w213), .x(w212) );
	dmg_not g41 (.a(w265), .x(w266) );
	dmg_not g42 (.a(w151), .x(w319) );
	dmg_not g43 (.a(w243), .x(w156) );
	dmg_not g44 (.a(w309), .x(w308) );
	dmg_not g45 (.a(w274), .x(w130) );
	dmg_not g46 (.a(w215), .x(w273) );
	dmg_not g47 (.a(w203), .x(w204) );
	dmg_not g48 (.a(w205), .x(w271) );
	dmg_not g49 (.a(w63), .x(w29) );
	dmg_not g50 (.a(w16), .x(w12) );
	dmg_not g51 (.a(w235), .x(w234) );
	dmg_not g52 (.a(w10), .x(w9) );
	dmg_nor g53 (.a(w36), .b(w2), .x(w1) );
	dmg_nor g54 (.a(w36), .b(w365), .x(w292) );
	dmg_nor g55 (.a(w36), .b(w230), .x(w291) );
	dmg_nor g56 (.a(w260), .b(w36), .x(w346) );
	dmg_nor g57 (.a(w242), .b(w277), .x(w278) );
	dmg_nor g58 (.a(w279), .b(w187), .x(w186) );
	dmg_nor g59 (.a(w29), .b(w356), .x(w15) );
	dmg_nor g60 (.a(w29), .b(w232), .x(w233) );
	dmg_nor g61 (.a(w29), .b(w18), .x(w17) );
	dmg_nor g62 (.a(w29), .b(w91), .x(w92) );
	dmg_nor g63 (.a(w29), .b(w335), .x(w334) );
	dmg_nor g64 (.a(w36), .b(w288), .x(w289) );
	dmg_nor g65 (.a(w89), .b(w43), .x(w42) );
	dmg_nor g66 (.a(w36), .b(w196), .x(w216) );
	dmg_nor g67 (.a(w36), .b(w42), .x(w41) );
	dmg_nor g68 (.a(w133), .b(w127), .x(w126) );
	dmg_nor g69 (.a(w36), .b(w26), .x(w268) );
	dmg_nor g70 (.a(w29), .b(w122), .x(w351) );
	dmg_nor g71 (.a(w29), .b(w121), .x(w350) );
	dmg_nor g72 (.a(w29), .b(w30), .x(w328) );
	dmg_nor g73 (.a(w263), .b(w215), .x(w198) );
	dmg_nor g74 (.a(w14), .b(w13), .x(w357) );
	dmg_nor g75 (.a(w36), .b(w227), .x(w270) );
	dmg_nor g76 (.a(w36), .b(w237), .x(w294) );
	dmg_nand g77 (.a(w2), .b(w8), .x(w7) );
	dmg_nand g78 (.a(w365), .b(w8), .x(w290) );
	dmg_nand g79 (.a(w230), .b(w8), .x(w51) );
	dmg_nand g80 (.a(w36), .b(w261), .x(w302) );
	dmg_nand g81 (.a(w321), .b(w322), .x(w183) );
	dmg_nand g82 (.a(w322), .b(w188), .x(w285) );
	dmg_nand g83 (.a(w196), .b(w8), .x(w40) );
	dmg_nand g84 (.a(w42), .b(w8), .x(w35) );
	dmg_nand g85 (.a(w26), .b(w8), .x(w267) );
	dmg_nand g86 (.a(w311), .b(w184), .x(w181) );
	dmg_nand g87 (.a(w185), .b(w284), .x(w283) );
	dmg_nand g88 (.a(w185), .b(w190), .x(w170) );
	dmg_nand g89 (.a(w227), .b(w8), .x(w236) );
	dmg_nand g90 (.a(w237), .b(w8), .x(w293) );
	dmg_bufif0 g91 (.a0(w50), .n_ena(w8), .a1(w50), .x(w49) );
	dmg_bufif0 g92 (.a0(w5), .n_ena(w8), .a1(w5), .x(w4) );
	dmg_bufif0 g93 (.a0(w234), .n_ena(w8), .a1(w234), .x(w272) );
	dmg_bufif0 g94 (.a0(w9), .n_ena(w8), .a1(w9), .x(w48) );
	dmg_bufif0 g95 (.a0(w11), .n_ena(w8), .a1(w11), .x(w229) );
	dmg_bufif0 g96 (.a0(w266), .n_ena(w8), .a1(w266), .x(w28) );
	dmg_latch g97 (.ena(w130), .d(w49), .q(w209) );
	dmg_latch g98 (.ena(w130), .d(w48), .q(w208) );
	dmg_latch g99 (.ena(w130), .d(w272), .q(w238) );
	dmg_latch g100 (.ena(w130), .d(w4), .q(w3) );
	dmg_latch g101 (.ena(w130), .d(w229), .q(w228) );
	dmg_latch g102 (.ena(w151), .d(w131), .nq(w154) );
	dmg_latch g103 (.ena(w151), .d(w162), .nq(w165) );
	dmg_latch g104 (.ena(w130), .d(w28), .q(w27) );
	dmg_latch g105 (.ena(w151), .d(w152), .nq(w353) );
	dmg_latch g106 (.ena(w151), .d(w164), .nq(w318) );
	dmg_latch g107 (.ena(w130), .d(w320), .q(w339) );
	dmg_latch g108 (.ena(w151), .d(w153), .nq(w326) );
	dmg_bufif0 g109 (.a0(w212), .n_ena(w8), .a1(w212), .x(w320) );
	dmg_dffr g110 (.clk(w74), .nr1(w12), .d(w14), .nr2(w12), .nq(w13) );
	dmg_dffr g111 (.clk(w225), .nr1(w63), .d(w68), .nr2(w63), .nq(w338), .q(w337) );
	dmg_dffr g112 (.clk(w360), .nr1(w177), .d(w171), .nr2(w177), .nq(w171), .q(w172) );
	dmg_dffr g113 (.clk(w367), .nr1(w177), .d(w176), .nr2(w177), .nq(w176), .q(w175) );
	dmg_dffr g114 (.clk(w340), .nr1(w177), .d(w246), .nr2(w177), .nq(w246), .q(w247) );
	dmg_dffr g115 (.clk(w361), .nr1(w177), .d(w280), .nr2(w177), .nq(w280), .q(w174) );
	dmg_dffr g116 (.clk(w279), .nr1(w188), .d(w278), .nr2(w188), .q(w366) );
	dmg_dffr g117 (.clk(w323), .nr1(w188), .d(w366), .nr2(w188), .nq(w322) );
	dmg_dffr g118 (.clk(w80), .nr1(w76), .d(w77), .nr2(w76), .nq(w77), .q(w314) );
	dmg_dffr g119 (.clk(w104), .nr1(w76), .d(w80), .nr2(w76), .nq(w80), .q(w79) );
	dmg_dffr g120 (.clk(w77), .nr1(w76), .d(w316), .nr2(w76), .nq(w316), .q(w315) );
	dmg_dffr g121 (.clk(w316), .nr1(w76), .d(w115), .nr2(w76), .nq(w115), .q(w114) );
	dmg_dffr g122 (.clk(w218), .nr1(w76), .d(w142), .nr2(w76), .nq(w142), .q(w143) );
	dmg_dffr g123 (.clk(w195), .nr1(w76), .d(w75), .nr2(w76), .nq(w75), .q(w219) );
	dmg_dffr g124 (.clk(w225), .nr1(w63), .d(w95), .nr2(w63), .nq(w97), .q(w96) );
	dmg_dffr g125 (.clk(w223), .nr1(w61), .d(w62), .nr2(w61), .nq(w62), .q(w141) );
	dmg_dffr g126 (.clk(w225), .nr1(w63), .d(w23), .nr2(w63), .nq(w331), .q(w224) );
	dmg_dffr g127 (.clk(w330), .nr1(w61), .d(w60), .nr2(w61), .nq(w60), .q(w59) );
	dmg_dffr g128 (.clk(w62), .nr1(w61), .d(w330), .nr2(w61), .nq(w330) );
	dmg_dffr g129 (.clk(w142), .nr1(w76), .d(w195), .nr2(w76), .nq(w195) );
	dmg_dffr g130 (.clk(w37), .nr1(w76), .d(w218), .nr2(w76), .nq(w218) );
	dmg_dffr g131 (.clk(w74), .nr1(w76), .d(w354), .nr2(w76), .nq(w354) );
	dmg_dffr g132 (.clk(w354), .nr1(w76), .d(w37), .nr2(w76), .nq(w37), .q(w81) );
	dmg_dffr g133 (.clk(w88), .nr1(w76), .d(w104), .nr2(w76), .nq(w104), .q(w105) );
	dmg_dffr g134 (.clk(w149), .nr1(w63), .d(w71), .nr2(w63), .nq(w127) );
	dmg_dffr g135 (.clk(w149), .nr1(w63), .d(w31), .nr2(w63), .nq(w347), .q(w83) );
	dmg_dffr g136 (.clk(w149), .nr1(w63), .d(w68), .nr2(w63), .nq(w253), .q(w252) );
	dmg_dffr g137 (.clk(w115), .nr1(w76), .d(w226), .nr2(w76), .nq(w226), .q(w137) );
	dmg_dffr g138 (.clk(w226), .nr1(w76), .d(w223), .nr2(w76), .nq(w223), .q(w116) );
	dmg_dffr g139 (.clk(w225), .nr1(w63), .d(w155), .nr2(w63), .nq(w303), .q(w363) );
	dmg_dffr g140 (.clk(w225), .nr1(w63), .d(w31), .nr2(w63), .nq(w222), .q(w336) );
	dmg_dffr g141 (.clk(w225), .nr1(w63), .d(w19), .nr2(w63), .nq(w98), .q(w99) );
	dmg_dffr g142 (.clk(w225), .nr1(w63), .d(w118), .nr2(w63), .nq(w119), .q(w120) );
	dmg_dffr g143 (.clk(w176), .nr1(w177), .d(w360), .nr2(w177), .nq(w360), .q(w281) );
	dmg_dffr g144 (.clk(w280), .nr1(w177), .d(w340), .nr2(w177), .nq(w340), .q(w173) );
	dmg_dffr g145 (.clk(w180), .nr1(w188), .d(w184), .nr2(w188), .q(w187) );
	dmg_dffr g146 (.clk(w279), .nr1(w188), .d(w183), .nr2(w188), .q(w185) );
	dmg_dffr g147 (.clk(w323), .nr1(w177), .d(w342), .nr2(w177), .nq(w189) );
	dmg_dffr g148 (.clk(w246), .nr1(w177), .d(w367), .nr2(w177), .nq(w367), .q(w343) );
	dmg_dffr g149 (.clk(w171), .nr1(w177), .d(w178), .nr2(w177), .nq(w178), .q(w179) );
	dmg_dffr g150 (.clk(w225), .nr1(w63), .d(w71), .nr2(w63), .nq(w297), .q(w298) );
	dmg_dffr g151 (.clk(w74), .nr1(w63), .d(w357), .nr2(w63), .q(w205) );
	dmg_dffsr g152 (.nset1(w301), .clk(w65), .nres(w64), .q(w164), .nset2(w301), .d(w21) );
	dmg_dffsr g153 (.nset1(w245), .clk(w259), .nres(w258), .q(w152), .nset2(w245), .d(w21) );
	dmg_dffsr g154 (.nset1(w255), .clk(w205), .nres(w352), .q(w153), .nset2(w255), .d(w21) );
	dmg_dffsr g155 (.nset1(w22), .clk(w358), .nres(w194), .q(w162), .nset2(w22), .d(w21) );
	dmg_dffsr g156 (.nset1(w134), .clk(w86), .nres(w135), .q(w131), .nset2(w134), .d(w21) );
	dmg_latchnq_comp g157 (.n_ena(w243), .d(w95), .ena(w156), .q(w158), .nq(w157) );
	dmg_latchnq_comp g158 (.n_ena(w243), .d(w23), .ena(w156), .q(w207), .nq(w355) );
	dmg_latchnq_comp g159 (.n_ena(w243), .d(w31), .ena(w156), .q(w239), .nq(w349) );
	dmg_latchnq_comp g160 (.n_ena(w243), .d(w118), .ena(w156), .q(w327), .nq(w348) );
	dmg_latchnq_comp g161 (.n_ena(w243), .d(w19), .ena(w156), .q(w211), .nq(w254) );
	dmg_latchnq_comp g162 (.n_ena(w243), .d(w68), .ena(w156), .q(w276), .nq(w129) );
	dmg_latchnq_comp g163 (.n_ena(w243), .d(w71), .ena(w156), .q(w282), .nq(w307) );
	dmg_latchnq_comp g164 (.n_ena(w243), .d(w155), .ena(w156), .q(w192), .nq(w244) );
	dmg_aon g165 (.a0(w273), .a1(w263), .b(w215), .x(w275) );
	dmg_aon g166 (.a0(w47), .a1(w325), .b(w201), .x(w200) );
	dmg_cnt g167 (.q(w14), .d(w350), .load(w16), .clk(w124), .nq(w123) );
	dmg_cnt g168 (.q(w125), .d(w328), .load(w16), .clk(w126), .nq(w220) );
	dmg_cnt g169 (.q(w333), .d(w334), .load(w16), .clk(w93), .nq(w94) );
	dmg_cnt g170 (.q(w329), .d(w17), .load(w16), .clk(w333), .nq(w332) );
	dmg_cnt g171 (.q(w93), .d(w92), .load(w16), .clk(w25), .nq(w24) );
	dmg_cnt g172 (.q(w124), .d(w351), .load(w16), .clk(w329), .nq(w231) );
	dmg_cnt g173 (.q(w73), .d(w15), .load(w16), .clk(w125), .nq(w296) );
	dmg_cnt g174 (.q(w25), .d(w233), .load(w16), .clk(w73), .nq(w72) );
	dmg_nor_latch g175 (.s(w242), .r(w285), .nq(w277) );
	dmg_nor_latch g176 (.s(w264), .r(w57), .nq(w58) );
	dmg_muxi g177 (.sel(w100), .d1(w298), .d0(w71), .q(w232) );
	dmg_muxi g178 (.sel(w100), .d1(w363), .d0(w155), .q(w121) );
	dmg_muxi g179 (.sel(w100), .d1(w120), .d0(w118), .q(w122) );
	dmg_muxi g180 (.sel(w100), .d1(w336), .d0(w31), .q(w30) );
	dmg_muxi g181 (.sel(w252), .d1(w84), .d0(w85), .q(w133) );
	dmg_muxi g182 (.sel(w83), .d1(w82), .d0(w78), .q(w85) );
	dmg_muxi g183 (.sel(w83), .d1(w53), .d0(w144), .q(w84) );
	dmg_muxi g184 (.sel(w36), .d1(w160), .d0(w47), .q(w46) );
	dmg_muxi g185 (.sel(w36), .d1(w217), .d0(w203), .q(w159) );
	dmg_muxi g186 (.sel(w100), .d1(w99), .d0(w19), .q(w18) );
	dmg_muxi g187 (.sel(w100), .d1(w224), .d0(w23), .q(w91) );
	dmg_muxi g188 (.sel(w100), .d1(w96), .d0(w95), .q(w335) );
	dmg_muxi g189 (.sel(w100), .d1(w337), .d0(w68), .q(w356) );
	dmg_and g190 (.a(w241), .b(w240), .x(w242) );
	dmg_and g191 (.a(w52), .b(w38), .x(w36) );
	dmg_and g192 (.a(w39), .b(w161), .x(w215) );
	dmg_and g193 (.a(w58), .b(w59), .x(w214) );
	dmg_and g194 (.a(w185), .b(w186), .x(w344) );
	dmg_and g195 (.a(w279), .b(w183), .x(w361) );
	dmg_and g196 (.a(w240), .b(w311), .x(w310) );
	dmg_not2 g197 (.a(w181), .x(w182) );
	dmg_not2 g198 (.a(w279), .x(w323) );
	dmg_not2 g199 (.a(w312), .x(w279) );
	dmg_not g200 (.a(w108), .x(w109) );
	dmg_not g201 (.a(w112), .x(w111) );
	dmg_not3 g202 (.a(w159), .x(w110) );
	dmg_not3 g203 (.a(w46), .x(w45) );
	dmg_and3 g204 (.a(w136), .b(w70), .c(w63), .x(w135) );
	dmg_and4 g205 (.a(w101), .b(w45), .c(w109), .d(w112), .x(w33) );
	dmg_and4 g206 (.a(w101), .b(w45), .c(w108), .d(w111), .x(w90) );
	dmg_and4 g207 (.a(w101), .b(w110), .c(w109), .d(w111), .x(w362) );
	dmg_and4 g208 (.a(w101), .b(w45), .c(w109), .d(w111), .x(w139) );
	dmg_and3 g209 (.a(w166), .b(w167), .c(w63), .x(w194) );
	dmg_and3 g210 (.a(w36), .b(w215), .c(w214), .x(w364) );
	dmg_and4 g211 (.a(w147), .b(w45), .c(w108), .d(w111), .x(w146) );
	dmg_and4 g212 (.a(w147), .b(w45), .c(w109), .d(w112), .x(w145) );
	dmg_notif1 g213 (.ena(w139), .a(w106), .x(w31) );
	dmg_notif1 g214 (.ena(w139), .a(w313), .x(w71) );
	dmg_notif1 g215 (.ena(w139), .a(w345), .x(w23) );
	dmg_notif1 g216 (.ena(w139), .a(w78), .x(w68) );
	dmg_notif1 g217 (.ena(w139), .a(w140), .x(w155) );
	dmg_notif1 g218 (.ena(w33), .a(w72), .x(w71) );
	dmg_notif1 g219 (.ena(w33), .a(w296), .x(w68) );
	dmg_notif1 g220 (.ena(w33), .a(w231), .x(w118) );
	dmg_notif1 g221 (.ena(w90), .a(w119), .x(w118) );
	dmg_notif1 g222 (.ena(w319), .a(w326), .x(w71) );
	dmg_notif1 g223 (.ena(w308), .a(w348), .x(w118) );
	dmg_notif1 g224 (.ena(w308), .a(w254), .x(w19) );
	dmg_notif1 g225 (.ena(w128), .a(w253), .x(w68) );
	dmg_notif1 g226 (.ena(w308), .a(w129), .x(w68) );
	dmg_notif1 g227 (.ena(w128), .a(w347), .x(w31) );
	dmg_notif1 g228 (.ena(w346), .a(w20), .x(w155) );
	dmg_notif1 g229 (.ena(w346), .a(w20), .x(w19) );
	dmg_notif1 g230 (.ena(w346), .a(w20), .x(w118) );
	dmg_notif1 g231 (.ena(w346), .a(w20), .x(w68) );
	dmg_notif1 g232 (.ena(w346), .a(w20), .x(w23) );
	dmg_notif1 g233 (.ena(w346), .a(w20), .x(w71) );
	dmg_notif1 g234 (.ena(w101), .a(w20), .x(w95) );
	dmg_notif1 g235 (.ena(w101), .a(w20), .x(w31) );
	dmg_notif1 g236 (.ena(w308), .a(w307), .x(w71) );
	dmg_notif1 g237 (.ena(w308), .a(w244), .x(w155) );
	dmg_notif1 g238 (.ena(w319), .a(w318), .x(w31) );
	dmg_notif1 g239 (.ena(w319), .a(w353), .x(w68) );
	dmg_notif1 g240 (.ena(w90), .a(w297), .x(w71) );
	dmg_notif1 g241 (.ena(w33), .a(w123), .x(w155) );
	dmg_notif1 g242 (.ena(w90), .a(w338), .x(w68) );
	dmg_notif1 g243 (.ena(w319), .a(w165), .x(w23) );
	dmg_notif1 g244 (.ena(w319), .a(w154), .x(w95) );
	dmg_notif1 g245 (.ena(w308), .a(w349), .x(w31) );
	dmg_notif1 g246 (.ena(w308), .a(w355), .x(w23) );
	dmg_notif1 g247 (.ena(w308), .a(w157), .x(w95) );
	dmg_notif1 g248 (.ena(w128), .a(w127), .x(w71) );
	dmg_notif1 g249 (.ena(w139), .a(w138), .x(w19) );
	dmg_notif1 g250 (.ena(w139), .a(w117), .x(w118) );
	dmg_notif1 g251 (.ena(w90), .a(w303), .x(w155) );
	dmg_notif1 g252 (.ena(w33), .a(w220), .x(w31) );
	dmg_notif1 g253 (.ena(w90), .a(w222), .x(w31) );
	dmg_notif1 g254 (.ena(w33), .a(w94), .x(w95) );
	dmg_notif1 g255 (.ena(w90), .a(w97), .x(w95) );
	dmg_notif1 g256 (.ena(w90), .a(w98), .x(w19) );
	dmg_notif1 g257 (.ena(w33), .a(w332), .x(w19) );
	dmg_notif1 g258 (.ena(w90), .a(w331), .x(w23) );
	dmg_notif1 g259 (.ena(w33), .a(w24), .x(w23) );
	dmg_notif1 g260 (.ena(w139), .a(w113), .x(w95) );
	dmg_nand6 g261 (.a(w174), .b(w173), .c(w247), .d(w343), .e(w175), .f(w179), .x(w341) );
	dmg_nand4 g262 (.a(w102), .b(w248), .c(w148), .d(w45), .x(w151) );
	dmg_nand4 g263 (.a(w102), .b(w248), .c(w148), .d(w110), .x(w150) );
	dmg_mux g264 (.sel(w36), .d1(w44), .d0(w43), .q(w261) );
	dmg_mux g265 (.sel(w87), .d1(w74), .d0(w75), .q(w88) );
	dmg_mux g266 (.sel(w89), .d1(w282), .d0(w339), .q(w288) );
	dmg_mux g267 (.sel(w89), .d1(w327), .d0(w27), .q(w26) );
	dmg_mux g268 (.sel(w89), .d1(w158), .d0(w209), .q(w230) );
	dmg_mux g269 (.sel(w89), .d1(w207), .d0(w208), .q(w365) );
	dmg_mux g270 (.sel(w89), .d1(w239), .d0(w238), .q(w237) );
	dmg_mux g271 (.sel(w89), .d1(w211), .d0(w3), .q(w2) );
	dmg_mux g272 (.sel(w89), .d1(w276), .d0(w228), .q(w227) );
	dmg_nand3 g273 (.a(w183), .b(w189), .c(w188), .x(w321) );
	dmg_nand3 g274 (.a(w47), .b(w263), .c(w206), .x(w262) );
	dmg_and3 g275 (.a(w300), .b(w193), .c(w63), .x(w64) );
	dmg_or g276 (.a(w204), .b(w198), .x(w197) );
	dmg_or g277 (.a(w68), .b(w32), .x(w67) );
	dmg_and3 g278 (.a(w306), .b(w304), .c(w148), .x(w101) );
	dmg_nand g279 (.a(w288), .b(w8), .x(w34) );
	dmg_or g280 (.a(w71), .b(w32), .x(w221) );
	dmg_nand3 g281 (.a(w69), .b(w167), .c(w23), .x(w22) );
	dmg_nand4 g282 (.a(w112), .b(w109), .c(w110), .d(w101), .x(w100) );
	dmg_nand4 g283 (.a(w111), .b(w108), .c(w110), .d(w101), .x(w225) );
	dmg_nand3 g284 (.a(w69), .b(w70), .c(w95), .x(w134) );
	dmg_nand3 g285 (.a(w38), .b(w161), .c(w55), .x(w54) );
	dmg_const g286 (.q0(w20), .q1(w21) );
	dmg_nand3 g287 (.a(w69), .b(w66), .c(w68), .x(w245) );
	dmg_nand3 g288 (.a(w69), .b(w193), .c(w31), .x(w301) );
	dmg_nand3 g289 (.a(w210), .b(w63), .c(w271), .x(w16) );
	dmg_or g290 (.a(w206), .b(w100), .x(w210) );
	dmg_or g291 (.a(w198), .b(w199), .x(w43) );
	dmg_or g292 (.a(w31), .b(w32), .x(w300) );
	dmg_or g293 (.a(w197), .b(w89), .x(w196) );
	dmg_or g294 (.a(w23), .b(w32), .x(w166) );
	dmg_or g295 (.a(w95), .b(w150), .x(w136) );
	dmg_or g296 (.a(w55), .b(w56), .x(w57) );
	dmg_nor5 g297 (.a(w251), .b(w250), .c(w107), .d(w103), .e(w249), .x(w304) );
	dmg_nor4 g298 (.a(w251), .b(w250), .c(w107), .d(w103), .x(w102) );
	dmg_and3 g299 (.a(w305), .b(w304), .c(w148), .x(w147) );
	dmg_and4 g300 (.a(w112), .b(w108), .c(w306), .d(w249), .x(w248) );
	dmg_and4 g301 (.a(w101), .b(w45), .c(w108), .d(w112), .x(w128) );
	dmg_nand4 g302 (.a(w112), .b(w108), .c(w110), .d(w101), .x(w149) );
	dmg_nand3 g303 (.a(w69), .b(w256), .c(w71), .x(w255) );
	dmg_and3 g304 (.a(w221), .b(w256), .c(w63), .x(w352) );
	dmg_nor3 g305 (.a(w211), .b(w327), .c(w191), .x(w190) );
	dmg_and3 g306 (.a(w67), .b(w66), .c(w63), .x(w258) );
	dmg_nand4 g307 (.a(w112), .b(w109), .c(w110), .d(w147), .x(w359) );
	dmg_nand4 g308 (.a(w111), .b(w108), .c(w110), .d(w147), .x(w317) );
	dmg_nor3 g309 (.a(w56), .b(w55), .c(w362), .x(w76) );
endmodule // MMIO