module Arbiter (  clk2, n_reset2, cpu_mreq, ext_cs_en, cpu_wr_sync, a[0], a[1], d[7], d[6], d[5], d[4], d[3], d[2], d[1], d[0], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], cpu_wr, mmio_sel, boot_sel, n_DRV_HIGH_a[15], n_INPUT_a[15], DRV_LOW_a[15], n_cs_topad, CONST0, n_DRV_HIGH_nmwr, n_mwr, DRV_LOW_nmwr, n_DRV_HIGH_nmrd, n_mrd, DRV_LOW_nmrd, n_DRV_HIGH_nmcs, n_mcs, DRV_LOW_nmcs, n_DRV_HIGH_md[7], n_md_frompad[7], DRV_LOW_md[7], n_md_ena_pu, n_DRV_HIGH_md[6], n_md_frompad[6], DRV_LOW_md[6], n_DRV_HIGH_md[5], n_md_frompad[5], DRV_LOW_md[5], n_DRV_HIGH_md[4], n_md_frompad[4], DRV_LOW_md[4], n_DRV_HIGH_md[3], n_md_frompad[3], DRV_LOW_md[3], n_DRV_HIGH_md[2], n_md_frompad[2], DRV_LOW_md[2], n_DRV_HIGH_md[1], n_md_frompad[1], DRV_LOW_md[1], n_DRV_HIGH_md[0], DRV_LOW_md[0], n_md_frompad[0], n_DRV_HIGH_d[7], n_db_frompad[7], DRV_LOW_d[7], n_ena_pu_db, n_DRV_HIGH_d[6], n_db_frompad[6], DRV_LOW_d[6], n_DRV_HIGH_d[5], n_db_frompad[5], DRV_LOW_d[5], n_DRV_HIGH_d[4], n_db_frompad[4], DRV_LOW_d[4], n_DRV_HIGH_d[3], n_db_frompad[3], DRV_LOW_d[3], n_DRV_HIGH_d[2], n_db_frompad[2], DRV_LOW_d[2], n_DRV_HIGH_d[1], n_db_frompad[1], DRV_LOW_d[1], n_DRV_HIGH_d[0], n_db_frompad[0], DRV_LOW_d[0], soc_wr, soc_rd, vram_to_oam, dma_a[15], non_vram_mreq, test_1, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, ffxx, n_ppu_hard_reset, ppu_mode3, md[2], md[5], md[1], md[7], md[0], md[6], md[3], md[4], arb_unk1, arb_unk2, arb_unk3, from_ppu2_unk2, arb_unk4, arb_unk5, from_mmio_unk1, arb_SUGY, arb_SYZO, sp_bp_cys, tm_bp_cys, from_ppu1_RAWA, n_tm_bp_cys, arb_RYCU, cpu_vram_oam_rd, arb_SERA);

	input wire clk2;
	input wire n_reset2;
	input wire cpu_mreq;
	input wire ext_cs_en;
	input wire cpu_wr_sync;
	input wire a[0];
	input wire a[1];
	inout wire d[7];
	inout wire d[6];
	inout wire d[5];
	inout wire d[4];
	inout wire d[3];
	inout wire d[2];
	inout wire d[1];
	inout wire d[0];
	input wire a[2];
	input wire a[3];
	input wire a[4];
	input wire a[5];
	input wire a[6];
	input wire a[7];
	input wire a[8];
	input wire a[9];
	input wire a[10];
	input wire a[11];
	input wire a[12];
	input wire a[13];
	input wire a[14];
	input wire a[15];
	input wire cpu_wr;
	output wire mmio_sel;
	output wire boot_sel;
	output wire n_DRV_HIGH_a[15];
	input wire n_INPUT_a[15];
	output wire DRV_LOW_a[15];
	output wire n_cs_topad;
	output wire CONST0;
	output wire n_DRV_HIGH_nmwr;
	input wire n_mwr;
	output wire DRV_LOW_nmwr;
	output wire n_DRV_HIGH_nmrd;
	input wire n_mrd;
	output wire DRV_LOW_nmrd;
	output wire n_DRV_HIGH_nmcs;
	input wire n_mcs;
	output wire DRV_LOW_nmcs;
	output wire n_DRV_HIGH_md[7];
	input wire n_md_frompad[7];
	output wire DRV_LOW_md[7];
	output wire n_md_ena_pu;
	output wire n_DRV_HIGH_md[6];
	input wire n_md_frompad[6];
	output wire DRV_LOW_md[6];
	output wire n_DRV_HIGH_md[5];
	input wire n_md_frompad[5];
	output wire DRV_LOW_md[5];
	output wire n_DRV_HIGH_md[4];
	input wire n_md_frompad[4];
	output wire DRV_LOW_md[4];
	output wire n_DRV_HIGH_md[3];
	input wire n_md_frompad[3];
	output wire DRV_LOW_md[3];
	output wire n_DRV_HIGH_md[2];
	input wire n_md_frompad[2];
	output wire DRV_LOW_md[2];
	output wire n_DRV_HIGH_md[1];
	input wire n_md_frompad[1];
	output wire DRV_LOW_md[1];
	output wire n_DRV_HIGH_md[0];
	output wire DRV_LOW_md[0];
	input wire n_md_frompad[0];
	output wire n_DRV_HIGH_d[7];
	input wire n_db_frompad[7];
	output wire DRV_LOW_d[7];
	input wire n_ena_pu_db;
	output wire n_DRV_HIGH_d[6];
	input wire n_db_frompad[6];
	output wire DRV_LOW_d[6];
	output wire n_DRV_HIGH_d[5];
	input wire n_db_frompad[5];
	output wire DRV_LOW_d[5];
	output wire n_DRV_HIGH_d[4];
	input wire n_db_frompad[4];
	output wire DRV_LOW_d[4];
	output wire n_DRV_HIGH_d[3];
	input wire n_db_frompad[3];
	output wire DRV_LOW_d[3];
	output wire n_DRV_HIGH_d[2];
	input wire n_db_frompad[2];
	output wire DRV_LOW_d[2];
	output wire n_DRV_HIGH_d[1];
	input wire n_db_frompad[1];
	output wire DRV_LOW_d[1];
	output wire n_DRV_HIGH_d[0];
	input wire n_db_frompad[0];
	output wire DRV_LOW_d[0];
	input wire soc_wr;
	input wire soc_rd;
	input wire vram_to_oam;
	input wire dma_a[15];
	output wire non_vram_mreq;
	input wire test_1;
	input wire n_extdb_to_intdb;
	input wire n_dblatch_to_intdb;
	input wire n_intdb_to_extdb;
	output wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ppu_mode3;
	inout wire md[2];
	inout wire md[5];
	inout wire md[1];
	inout wire md[7];
	inout wire md[0];
	inout wire md[6];
	inout wire md[3];
	inout wire md[4];
	output wire arb_unk1;
	output wire arb_unk2;
	output wire arb_unk3;
	input wire from_ppu2_unk2;
	output wire arb_unk4;
	output wire arb_unk5;
	input wire from_mmio_unk1;
	output wire arb_SUGY;
	output wire arb_SYZO;
	input wire sp_bp_cys;
	input wire tm_bp_cys;
	input wire from_ppu1_RAWA;
	input wire n_tm_bp_cys;
	output wire arb_RYCU;
	input wire cpu_vram_oam_rd;
	output wire arb_SERA;

endmodule // Arbiter