module PPU1 (  a, d, n_ma, n_lcd_ld1, n_lcd_ld0, n_lcd_cpg, n_lcd_cp, n_lcd_st, n_lcd_cpl, n_lcd_fr, n_lcd_s, CONST0, n_dma_phi, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, ffxx, n_ppu_hard_reset, ff46, 
	nma, fexx, ff43, ff42, sprite_x_flip, sprite_x_match, bp_sel, ppu_mode3, 
	md, v, FF43_D1, FF43_D0, n_ppu_clk, FF43_D2, h, ppu_mode2, vbl, stop_oam_eval, obj_color, vclk2, h_restart, obj_prio_ck, obj_prio, n_ppu_reset, n_dma_phi2_latched, FF40_D3, FF40_D2, in_window, 
	FF40_D1, sp_bp_cys, tm_bp_cys, n_sp_bp_mrd, n_tm_bp_cys, arb_fexx_ffxx, ppu_int_stat, ppu_int_vbl, oam_mode3_bl_pch, bp_cy, tm_cy, oam_mode3_nrd, ppu1_ma0, oam_rd_ck, oam_xattr_latch_cck, oam_addr_ck);

	input wire [12:0] a;
	inout wire [7:0] d;
	output wire [12:0] n_ma;
	output wire n_lcd_ld1;
	output wire n_lcd_ld0;
	output wire n_lcd_cpg;
	output wire n_lcd_cp;
	output wire n_lcd_st;
	output wire n_lcd_cpl;
	output wire n_lcd_fr;
	output wire n_lcd_s;
	inout wire CONST0;
	input wire n_dma_phi;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire ppu_clk;
	input wire vram_to_oam;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	output wire ff46;
	inout wire [12:0] nma;
	output wire fexx;
	output wire ff43;
	output wire ff42;
	input wire sprite_x_flip;
	input wire sprite_x_match;
	output wire bp_sel;
	output wire ppu_mode3;
	inout wire [7:0] md;
	input wire FF43_D1;
	input wire FF43_D0;
	input wire n_ppu_clk;
	input wire FF43_D2;
	input wire ppu_mode2;
	output wire vbl;
	input wire stop_oam_eval;
	input wire obj_color;
	output wire vclk2;
	input wire obj_prio;
	output wire n_ppu_reset;
	output wire FF40_D3;
	output wire FF40_D2;
	output wire in_window;
	output wire FF40_D1;
	output wire sp_bp_cys;
	output wire tm_bp_cys;
	output wire n_tm_bp_cys;
	input wire arb_fexx_ffxx;
	output wire ppu_int_stat;
	output wire ppu_int_vbl;
	output wire bp_cy;
	output wire tm_cy;
	input wire h_restart;
	output wire obj_prio_ck;
	output wire n_dma_phi2_latched;
	output wire ppu1_ma0;
	output wire n_sp_bp_mrd; 		// to arb

	output wire oam_mode3_nrd;  		// is low when OAM is read during MODE3 (pixel transfer stage)
	output wire oam_mode3_bl_pch;
	// @msinger: I guess you already noticed yourself that XUJY(oam_mode3_bl_pch) is the same as XUJA(oam_mode3_nrd), but it is low for a little bit longer.
	// I don't know why it is longer, but it seems to be used to control the OAM bitline precharging during MODE3. It disables the precharging temporarily so that the read access can be performed.   (#328)

	// OAM Clocks
	output wire oam_rd_ck;
	output wire oam_xattr_latch_cck;
	output wire oam_addr_ck;

	// H/V

	output wire [7:0] h;
	output wire [7:0] v;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;
	wire w974;
	wire w975;
	wire w976;
	wire w977;
	wire w978;
	wire w979;
	wire w980;

	assign n_tm_bp_cys = w765;
	assign tm_bp_cys = w212;
	assign n_sp_bp_mrd = w552;
	assign md[5] = w311;
	assign md[2] = w121;
	assign md[1] = w553;
	assign md[7] = w120;
	assign w769 = arb_fexx_ffxx;
	assign md[6] = w554;
	assign md[3] = w218;
	assign w555 = a[12];
	assign w593 = a[11];
	assign w594 = a[9];
	assign w333 = a[8];
	assign md[0] = w332;
	assign w595 = a[10];
	assign sp_bp_cys = w123;
	assign ppu_int_vbl = w380;
	assign ppu_int_stat = w379;
	assign w574 = a[4];
	assign w575 = vram_to_oam;
	assign ff46 = w641;
	assign w128 = ffxx;
	assign w129 = a[3];
	assign w919 = a[0];
	assign w130 = a[1];
	assign nma[8] = w126;
	assign w127 = a[6];
	assign ppu_mode3 = w231;
	assign w134 = a[7];
	assign nma[7] = w135;
	assign w133 = a[5];
	assign w132 = a[2];
	assign nma[1] = w131;
	assign w136 = n_ppu_hard_reset;
	assign nma[9] = w566;
	assign fexx = w824;
	assign nma[0] = w272;
	assign ff43 = w850;
	assign nma[4] = w517;
	assign nma[12] = w65;
	assign nma[6] = w271;
	assign nma[5] = w49;
	assign ff42 = w270;
	assign nma[11] = w48;
	assign w59 = ppu_rd;
	assign nma[10] = w60;
	assign w152 = ppu_wr;
	assign w153 = sprite_x_flip;
	assign w853 = n_dma_phi;
	assign n_dma_phi2_latched = w74;
	assign nma[3] = w277;
	assign nma[2] = w154;
	assign w620 = sprite_x_match;
	assign oam_mode3_bl_pch = w224;
	assign bp_sel = w223;
	assign w825 = FF43_D1;
	assign v[7] = w77;
	assign bp_cy = w210;
	assign tm_cy = w211;
	assign w11 = FF43_D0;
	assign d[4] = w68;
	assign w319 = n_ppu_clk;
	assign d[7] = w79;
	assign w828 = FF43_D2;
	assign h[3] = w171;
	assign v[6] = w172;
	assign d[1] = w12;
	assign d[3] = w52;
	assign d[6] = w249;
	assign d[2] = w91;
	assign d[0] = w13;
	assign d[5] = w341;
	assign CONST0 = w14;
	assign v[4] = w281;
	assign v[0] = w252;
	assign h[4] = w814;
	assign h[6] = w375;
	assign h[7] = w624;
	assign FF40_D3 = w54;
	assign FF40_D2 = w55;
	assign in_window = w145;
	assign h[5] = w551;
	assign w851 = h_restart;
	assign oam_mode3_nrd = w339;
	assign v[3] = w255;
	assign ppu1_ma0 = w244;
	assign v[2] = w245;
	assign h[2] = w369;
	assign oam_rd_ck = w287;
	assign v[1] = w286;
	assign v[5] = w361;
	assign oam_xattr_latch_cck = w362;
	assign FF40_D1 = w829;
	assign oam_addr_ck = w496;
	assign h[0] = w497;
	assign w368 = ppu_mode2;
	assign h[1] = w521;
	assign vbl = w960;
	assign w533 = stop_oam_eval;
	assign w199 = obj_color;
	assign vclk2 = w687;
	assign w527 = obj_prio;
	assign obj_prio_ck = w293;
	assign n_ppu_reset = w148;
	assign w367 = ppu_clk;
	assign n_ma[11] = w584;
	assign n_ma[9] = w585;
	assign n_ma[8] = w796;
	assign n_lcd_cpl = w781;
	assign n_lcd_ld1 = w4;
	assign n_lcd_cp = w5;
	assign n_lcd_st = w531;
	assign n_lcd_ld0 = w530;
	assign n_lcd_cpg = w950;
	assign n_ma[10] = w62;
	assign n_ma[12] = w63;
	assign n_lcd_fr = w421;
	assign n_lcd_s = w422;
	assign n_ma[6] = w472;
	assign n_ma[5] = w51;
	assign n_ma[7] = w514;
	assign n_ma[3] = w279;
	assign n_ma[2] = w156;
	assign n_ma[4] = w471;
	assign n_ma[1] = w390;
	assign n_ma[0] = w802;
	assign md[4] = w217;

	// Instances

	dmg_not g1 (.a(w764), .x(w325) );
	dmg_not g2 (.a(w216), .x(w925) );
	dmg_not g3 (.a(w324), .x(w326) );
	dmg_not g4 (.a(w666), .x(w665) );
	dmg_not g5 (.a(w664), .x(w663) );
	dmg_not g6 (.a(w331), .x(w330) );
	dmg_not g7 (.a(w219), .x(w119) );
	dmg_not g8 (.a(w317), .x(w761) );
	dmg_not g9 (.a(w220), .x(w219) );
	dmg_not g10 (.a(w320), .x(w166) );
	dmg_not g11 (.a(w468), .x(w469) );
	dmg_not g12 (.a(w231), .x(w667) );
	dmg_not g13 (.a(w862), .x(w95) );
	dmg_not g14 (.a(w807), .x(w93) );
	dmg_not g15 (.a(w319), .x(w600) );
	dmg_not g16 (.a(w93), .x(w92) );
	dmg_not g17 (.a(w148), .x(w409) );
	dmg_not g18 (.a(w409), .x(w424) );
	dmg_not g19 (.a(w199), .x(w947) );
	dmg_not g20 (.a(w108), .x(w733) );
	dmg_not g21 (.a(w199), .x(w774) );
	dmg_not g22 (.a(w419), .x(w940) );
	dmg_not g23 (.a(w19), .x(w437) );
	dmg_not g24 (.a(w436), .x(w188) );
	dmg_not g25 (.a(w28), .x(w27) );
	dmg_not g26 (.a(w18), .x(w939) );
	dmg_not g27 (.a(w399), .x(w347) );
	dmg_not g28 (.a(w22), .x(w21) );
	dmg_not g29 (.a(w938), .x(w393) );
	dmg_not g30 (.a(w202), .x(w201) );
	dmg_not g31 (.a(w16), .x(w444) );
	dmg_not g32 (.a(w443), .x(w17) );
	dmg_not g33 (.a(w396), .x(w395) );
	dmg_not g34 (.a(w394), .x(w397) );
	dmg_not g35 (.a(w199), .x(w528) );
	dmg_not g36 (.a(w20), .x(w487) );
	dmg_not g37 (.a(w110), .x(w111) );
	dmg_not g38 (.a(w458), .x(w457) );
	dmg_not g39 (.a(w888), .x(w887) );
	dmg_not g40 (.a(w295), .x(w413) );
	dmg_not g41 (.a(w426), .x(w749) );
	dmg_not g42 (.a(w949), .x(w628) );
	dmg_not g43 (.a(w626), .x(w627) );
	dmg_not g44 (.a(w147), .x(w146) );
	dmg_not g45 (.a(w633), .x(w808) );
	dmg_not g46 (.a(w461), .x(w460) );
	dmg_not g47 (.a(w464), .x(w462) );
	dmg_not g48 (.a(w861), .x(w222) );
	dmg_not g49 (.a(w328), .x(w327) );
	dmg_not g50 (.a(w118), .x(w315) );
	dmg_not g51 (.a(w214), .x(w213) );
	dmg_not g52 (.a(w582), .x(w552) );
	dmg_not g53 (.a(w46), .x(w45) );
	dmg_not g54 (.a(w766), .x(w967) );
	dmg_not g55 (.a(w767), .x(w860) );
	dmg_not g56 (.a(w770), .x(w556) );
	dmg_not g57 (.a(w858), .x(w917) );
	dmg_not g58 (.a(w503), .x(w504) );
	dmg_not g59 (.a(w148), .x(w535) );
	dmg_not g60 (.a(w48), .x(w583) );
	dmg_not g61 (.a(w630), .x(w632) );
	dmg_not g62 (.a(w630), .x(w631) );
	dmg_not g63 (.a(w65), .x(w64) );
	dmg_not g64 (.a(w965), .x(w966) );
	dmg_not g65 (.a(w60), .x(w61) );
	dmg_not g66 (.a(w601), .x(w602) );
	dmg_not g67 (.a(w601), .x(w613) );
	dmg_not g68 (.a(w199), .x(w951) );
	dmg_not g69 (.a(w449), .x(w34) );
	dmg_not g70 (.a(w447), .x(w943) );
	dmg_not g71 (.a(w199), .x(w792) );
	dmg_not g72 (.a(w722), .x(w200) );
	dmg_not g73 (.a(w706), .x(w702) );
	dmg_not g74 (.a(w711), .x(w704) );
	dmg_not g75 (.a(w707), .x(w703) );
	dmg_not g76 (.a(w404), .x(w795) );
	dmg_not g77 (.a(w712), .x(w676) );
	dmg_not g78 (.a(w199), .x(w952) );
	dmg_not g79 (.a(w527), .x(w717) );
	dmg_not g80 (.a(w194), .x(w195) );
	dmg_not g81 (.a(w527), .x(w691) );
	dmg_not g82 (.a(w651), .x(w453) );
	dmg_not g83 (.a(w109), .x(w108) );
	dmg_not g84 (.a(w229), .x(w868) );
	dmg_not g85 (.a(w231), .x(w598) );
	dmg_not g86 (.a(w175), .x(w207) );
	dmg_not g87 (.a(w148), .x(w648) );
	dmg_not g88 (.a(w171), .x(w377) );
	dmg_not g89 (.a(w654), .x(w378) );
	dmg_not g90 (.a(w656), .x(w657) );
	dmg_not g91 (.a(w180), .x(w181) );
	dmg_not g92 (.a(w657), .x(w658) );
	dmg_not g93 (.a(w600), .x(w164) );
	dmg_not g94 (.a(w596), .x(w913) );
	dmg_not g95 (.a(w565), .x(w969) );
	dmg_not g96 (.a(w145), .x(w800) );
	dmg_not g97 (.a(w267), .x(w266) );
	dmg_not g98 (.a(w236), .x(w162) );
	dmg_not g99 (.a(w567), .x(w265) );
	dmg_not g100 (.a(w799), .x(w264) );
	dmg_not g101 (.a(w58), .x(w57) );
	dmg_not g102 (.a(w927), .x(w67) );
	dmg_not g103 (.a(w281), .x(w974) );
	dmg_not g104 (.a(w252), .x(w973) );
	dmg_not g105 (.a(w72), .x(w71) );
	dmg_not g106 (.a(w603), .x(w842) );
	dmg_not g107 (.a(w32), .x(w830) );
	dmg_not g108 (.a(w305), .x(w304) );
	dmg_not g109 (.a(w355), .x(w353) );
	dmg_not g110 (.a(w356), .x(w354) );
	dmg_not g111 (.a(w442), .x(w355) );
	dmg_not g112 (.a(w694), .x(w695) );
	dmg_not g113 (.a(w695), .x(w451) );
	dmg_not g114 (.a(w527), .x(w833) );
	dmg_not g115 (.a(w527), .x(w956) );
	dmg_not g116 (.a(w69), .x(w70) );
	dmg_not g117 (.a(w527), .x(w841) );
	dmg_not g118 (.a(w527), .x(w839) );
	dmg_not g119 (.a(w31), .x(w30) );
	dmg_not g120 (.a(w846), .x(w69) );
	dmg_not g121 (.a(w962), .x(w343) );
	dmg_not g122 (.a(w293), .x(w36) );
	dmg_not g123 (.a(w527), .x(w686) );
	dmg_not g124 (.a(w366), .x(w365) );
	dmg_not g125 (.a(w367), .x(w366) );
	dmg_not g126 (.a(w527), .x(w688) );
	dmg_not g127 (.a(w137), .x(w82) );
	dmg_not g128 (.a(w84), .x(w83) );
	dmg_not g129 (.a(w365), .x(w364) );
	dmg_not g130 (.a(w363), .x(w362) );
	dmg_not g131 (.a(w361), .x(w360) );
	dmg_not g132 (.a(w172), .x(w337) );
	dmg_not g133 (.a(w77), .x(w78) );
	dmg_not g134 (.a(w255), .x(w338) );
	dmg_not g135 (.a(w340), .x(w339) );
	dmg_not g136 (.a(w286), .x(w285) );
	dmg_not g137 (.a(w853), .x(w150) );
	dmg_not g138 (.a(w84), .x(w85) );
	dmg_not g139 (.a(w85), .x(w539) );
	dmg_not g140 (.a(w851), .x(w541) );
	dmg_not g141 (.a(w225), .x(w224) );
	dmg_not g142 (.a(w623), .x(w622) );
	dmg_not g143 (.a(w620), .x(w621) );
	dmg_not g144 (.a(w137), .x(w138) );
	dmg_not g145 (.a(w222), .x(w223) );
	dmg_not g146 (.a(w336), .x(w274) );
	dmg_not g147 (.a(w132), .x(w799) );
	dmg_not g148 (.a(w130), .x(w567) );
	dmg_not g149 (.a(w129), .x(w236) );
	dmg_not g150 (.a(w919), .x(w267) );
	dmg_not g151 (.a(w126), .x(w797) );
	dmg_not g152 (.a(w921), .x(w372) );
	dmg_not g153 (.a(w538), .x(w88) );
	dmg_not g154 (.a(w296), .x(w295) );
	dmg_not g155 (.a(w261), .x(w260) );
	dmg_not g156 (.a(w159), .x(w158) );
	dmg_not g157 (.a(w566), .x(w586) );
	dmg_not g158 (.a(w297), .x(w110) );
	dmg_not g159 (.a(w71), .x(w248) );
	dmg_not g160 (.a(w716), .x(w713) );
	dmg_not g161 (.a(w400), .x(w705) );
	dmg_not g162 (.a(w935), .x(w401) );
	dmg_not g163 (.a(w405), .x(w794) );
	dmg_not g164 (.a(w699), .x(w356) );
	dmg_not g165 (.a(w199), .x(w793) );
	dmg_not g166 (.a(w693), .x(w694) );
	dmg_not g167 (.a(w728), .x(w727) );
	dmg_not g168 (.a(w199), .x(w867) );
	dmg_not g169 (.a(w669), .x(w866) );
	dmg_not g170 (.a(w513), .x(w975) );
	dmg_not g171 (.a(w451), .x(w309) );
	dmg_not g172 (.a(w698), .x(w475) );
	dmg_not g173 (.a(w308), .x(w953) );
	dmg_not g174 (.a(w33), .x(w872) );
	dmg_not g175 (.a(w35), .x(w306) );
	dmg_not g176 (.a(w668), .x(w458) );
	dmg_not g177 (.a(w177), .x(w656) );
	dmg_not g178 (.a(w637), .x(w386) );
	dmg_not g179 (.a(w657), .x(w502) );
	dmg_not g180 (.a(w183), .x(w165) );
	dmg_not g181 (.a(w128), .x(w854) );
	dmg_not g182 (.a(w562), .x(w588) );
	dmg_not g183 (.a(w231), .x(w8) );
	dmg_not g184 (.a(w510), .x(w511) );
	dmg_not g185 (.a(w148), .x(w176) );
	dmg_not g186 (.a(w613), .x(w612) );
	dmg_not g187 (.a(w614), .x(w532) );
	dmg_not g188 (.a(w743), .x(w741) );
	dmg_not g189 (.a(w740), .x(w175) );
	dmg_not g190 (.a(w203), .x(w888) );
	dmg_not g191 (.a(w887), .x(w449) );
	dmg_not g192 (.a(w699), .x(w789) );
	dmg_not g193 (.a(w442), .x(w394) );
	dmg_not g194 (.a(w438), .x(w104) );
	dmg_not g195 (.a(w245), .x(w259) );
	dmg_not g196 (.a(w277), .x(w278) );
	dmg_not g197 (.a(w154), .x(w155) );
	dmg_not g198 (.a(w88), .x(w818) );
	dmg_not g199 (.a(w271), .x(w895) );
	dmg_not g200 (.a(w49), .x(w50) );
	dmg_not g201 (.a(w319), .x(w819) );
	dmg_not g202 (.a(w319), .x(w897) );
	dmg_not g203 (.a(w319), .x(w659) );
	dmg_not g204 (.a(w272), .x(w801) );
	dmg_not g205 (.a(w517), .x(w518) );
	dmg_not g206 (.a(w135), .x(w515) );
	dmg_not g207 (.a(w131), .x(w389) );
	dmg_not g208 (.a(w221), .x(w220) );
	dmg_not g209 (.a(w764), .x(w765) );
	dmg_dffsr g210 (.nset1(w805), .nset2(w805), .clk(w44), .nres(w937), .d(w25), .q(w721) );
	dmg_dffsr g211 (.nset1(w24), .nset2(w24), .clk(w44), .nres(w398), .d(w23), .q(w25) );
	dmg_dffsr g212 (.nset1(w29), .nset2(w29), .clk(w44), .nres(w977), .d(w473), .q(w28) );
	dmg_dffsr g213 (.nset1(w215), .nset2(w215), .clk(w44), .nres(w114), .d(w322), .q(w115) );
	dmg_dffsr g214 (.nset1(w117), .nset2(w117), .clk(w44), .nres(w758), .d(w116), .q(w757) );
	dmg_dffsr g215 (.nset1(w759), .nset2(w759), .clk(w44), .nres(w821), .d(w923), .q(w924) );
	dmg_dffsr g216 (.nset1(w196), .nset2(w196), .clk(w44), .nres(w777), .d(w197), .q(w776) );
	dmg_dffsr g217 (.nset1(w15), .nset2(w15), .clk(w44), .nres(w941), .d(w14), .q(w783) );
	dmg_dffsr g218 (.nset1(w942), .nset2(w942), .clk(w44), .nres(w787), .d(w14), .q(w784) );
	dmg_dffsr g219 (.nset1(w725), .nset2(w725), .clk(w44), .nres(w724), .d(w445), .q(w37) );
	dmg_dffsr g220 (.nset1(w674), .nset2(w674), .clk(w44), .nres(w790), .d(w673), .q(w729) );
	dmg_dffsr g221 (.nset1(w945), .nset2(w945), .clk(w44), .nres(w671), .d(w14), .q(w672) );
	dmg_dffsr g222 (.nset1(w590), .nset2(w590), .clk(w44), .nres(w768), .d(w589), .q(w859) );
	dmg_dffsr g223 (.nset1(w559), .nset2(w559), .clk(w44), .nres(w918), .d(w558), .q(w560) );
	dmg_dffsr g224 (.nset1(w910), .nset2(w910), .clk(w44), .nres(w911), .d(w909), .q(w563) );
	dmg_dffsr g225 (.nset1(w914), .nset2(w914), .clk(w44), .nres(w908), .d(w14), .q(w909) );
	dmg_dffsr g226 (.nset1(w680), .nset2(w680), .clk(w44), .nres(w681), .d(w679), .q(w682) );
	dmg_dffsr g227 (.nset1(w720), .nset2(w720), .clk(w44), .nres(w840), .d(w721), .q(w191) );
	dmg_dffsr g228 (.nset1(w928), .nset2(w928), .clk(w44), .nres(w934), .d(w190), .q(w930) );
	dmg_dffsr g229 (.nset1(w192), .nset2(w192), .clk(w44), .nres(w929), .d(w191), .q(w193) );
	dmg_dffsr g230 (.nset1(w844), .nset2(w844), .clk(w44), .nres(w845), .d(w39), .q(w40) );
	dmg_dffsr g231 (.nset1(w478), .nset2(w478), .clk(w44), .nres(w843), .d(w477), .q(w43) );
	dmg_dffsr g232 (.nset1(w303), .nset2(w303), .clk(w44), .nres(w685), .d(w684), .q(w302) );
	dmg_dffsr g233 (.nset1(w683), .nset2(w683), .clk(w44), .nres(w959), .d(w682), .q(w684) );
	dmg_dffsr g234 (.nset1(w677), .nset2(w677), .clk(w44), .nres(w715), .d(w38), .q(w39) );
	dmg_dffsr g235 (.nset1(w931), .nset2(w931), .clk(w44), .nres(w718), .d(w930), .q(w679) );
	dmg_dffsr g236 (.nset1(w955), .nset2(w955), .clk(w44), .nres(w476), .d(w193), .q(w477) );
	dmg_dffsr g237 (.nset1(w692), .nset2(w692), .clk(w44), .nres(w954), .d(w40), .q(w41) );
	dmg_dffsr g238 (.nset1(w870), .nset2(w870), .clk(w44), .nres(w871), .d(w41), .q(w42) );
	dmg_dffsr g239 (.nset1(w187), .nset2(w187), .clk(w44), .nres(w189), .d(w186), .q(w190) );
	dmg_dffsr g240 (.nset1(w301), .nset2(w301), .clk(w44), .nres(w690), .d(w302), .q(w300) );
	dmg_dffsr g241 (.nset1(w299), .nset2(w299), .clk(w44), .nres(w689), .d(w300), .q(w298) );
	dmg_dffsr g242 (.nset1(w581), .nset2(w581), .clk(w44), .nres(w557), .d(w592), .q(w558) );
	dmg_dffsr g243 (.nset1(w564), .nset2(w564), .clk(w44), .nres(w968), .d(w563), .q(w589) );
	dmg_dffsr g244 (.nset1(w561), .nset2(w561), .clk(w44), .nres(w141), .d(w560), .q(w140) );
	dmg_dffsr g245 (.nset1(w591), .nset2(w591), .clk(w44), .nres(w912), .d(w859), .q(w592) );
	dmg_dffsr g246 (.nset1(w710), .nset2(w710), .clk(w44), .nres(w709), .d(w672), .q(w673) );
	dmg_dffsr g247 (.nset1(w730), .nset2(w730), .clk(w44), .nres(w731), .d(w729), .q(w791) );
	dmg_dffsr g248 (.nset1(w726), .nset2(w726), .clk(w44), .nres(w723), .d(w37), .q(w38) );
	dmg_dffsr g249 (.nset1(w675), .nset2(w675), .clk(w44), .nres(w198), .d(w791), .q(w197) );
	dmg_dffsr g250 (.nset1(w782), .nset2(w782), .clk(w44), .nres(w446), .d(w783), .q(w445) );
	dmg_dffsr g251 (.nset1(w312), .nset2(w312), .clk(w44), .nres(w112), .d(w757), .q(w756) );
	dmg_dffsr g252 (.nset1(w323), .nset2(w323), .clk(w44), .nres(w762), .d(w321), .q(w322) );
	dmg_dffsr g253 (.nset1(w662), .nset2(w662), .clk(w44), .nres(w661), .d(w115), .q(w116) );
	dmg_dffsr g254 (.nset1(w316), .nset2(w316), .clk(w44), .nres(w760), .d(w924), .q(w321) );
	dmg_dffsr g255 (.nset1(w329), .nset2(w329), .clk(w44), .nres(w763), .d(w14), .q(w923) );
	dmg_dffsr g256 (.nset1(w474), .nset2(w474), .clk(w44), .nres(w775), .d(w776), .q(w473) );
	dmg_dffsr g257 (.nset1(w785), .nset2(w785), .clk(w44), .nres(w788), .d(w784), .q(w23) );
	dmg_dffr g258 (.clk(w659), .nr1(w143), .nr2(w143), .d(w166), .nq(w318) );
	dmg_dffr g259 (.clk(w467), .nr1(w143), .nr2(w143), .d(w466), .nq(w466), .q(w468) );
	dmg_dffr g260 (.clk(w319), .nr1(w231), .nr2(w231), .d(w468), .q(w470) );
	dmg_dffr g261 (.clk(w412), .nr1(w257), .nr2(w257), .d(w258), .nq(w258), .q(w245) );
	dmg_dffr g262 (.clk(w258), .nr1(w257), .nr2(w257), .d(w256), .nq(w256), .q(w255) );
	dmg_dffr g263 (.clk(w256), .nr1(w257), .nr2(w257), .d(w280), .nq(w280), .q(w281) );
	dmg_dffr g264 (.clk(w280), .nr1(w257), .nr2(w257), .d(w411), .nq(w411), .q(w361) );
	dmg_dffr g265 (.clk(w493), .nr1(w257), .nr2(w257), .d(w76), .nq(w76), .q(w77) );
	dmg_dffr g266 (.clk(w697), .nr1(w696), .nr2(w696), .d(w976), .nq(w976) );
	dmg_dffr g267 (.clk(w940), .nr1(w696), .nr2(w696), .d(w697), .nq(w697) );
	dmg_dffr g268 (.clk(w739), .nr1(w424), .nr2(w424), .d(w738), .nq(w738), .q(w963) );
	dmg_dffr g269 (.clk(w513), .nr1(w424), .nr2(w424), .d(w419), .nq(w173), .q(w174) );
	dmg_dffr g270 (.clk(w319), .nr1(w148), .nr2(w148), .d(w147), .nq(w634) );
	dmg_dffr g271 (.clk(w819), .nr1(w231), .nr2(w231), .d(w810), .nq(w809) );
	dmg_dffr g272 (.clk(w897), .nr1(w148), .nr2(w148), .d(w168), .q(w536) );
	dmg_dffr g273 (.clk(w319), .nr1(w167), .nr2(w167), .d(w166), .q(w875) );
	dmg_dffr g274 (.clk(w465), .nr1(w143), .nr2(w143), .d(w922), .nq(w922), .q(w861) );
	dmg_dffr g275 (.clk(w319), .nr1(w231), .nr2(w231), .d(w755), .q(w907) );
	dmg_dffr g276 (.clk(w630), .nr1(w231), .nr2(w231), .d(w629), .nq(w916), .q(w755) );
	dmg_dffr g277 (.clk(w885), .nr1(w505), .nr2(w505), .d(w902), .nq(w902), .q(w883) );
	dmg_dffr g278 (.clk(w509), .nr1(w505), .nr2(w505), .d(w885), .nq(w885), .q(w884) );
	dmg_dffr g279 (.clk(w506), .nr1(w505), .nr2(w505), .d(w509), .nq(w509), .q(w508) );
	dmg_dffr g280 (.clk(w513), .nr1(w247), .nr2(w247), .d(w741), .q(w550) );
	dmg_dffr g281 (.clk(w975), .nr1(w424), .nr2(w424), .d(w732), .q(w419) );
	dmg_dffr g282 (.clk(w407), .nr1(w408), .nr2(w408), .d(w708), .nq(w708), .q(w935) );
	dmg_dffr g283 (.clk(w933), .nr1(w408), .nr2(w408), .d(w678), .nq(w678), .q(w707) );
	dmg_dffr g284 (.clk(w678), .nr1(w408), .nr2(w408), .d(w719), .nq(w719), .q(w711) );
	dmg_dffr g285 (.clk(w932), .nr1(w408), .nr2(w408), .d(w406), .nq(w406), .q(w405) );
	dmg_dffr g286 (.clk(w600), .nr1(w186), .nr2(w186), .d(w229), .nq(w240), .q(w205) );
	dmg_dffr g287 (.clk(w822), .nr1(w823), .nr2(w823), .d(w228), .nq(w228), .q(w229) );
	dmg_dffr g288 (.clk(w228), .nr1(w823), .nr2(w823), .d(w971), .nq(w971), .q(w526) );
	dmg_dffr g289 (.clk(w971), .nr1(w823), .nr2(w823), .d(w972), .nq(w972), .q(w227) );
	dmg_dffr g290 (.clk(w377), .nr1(w499), .nr2(w499), .d(w901), .q(w551) );
	dmg_dffr g291 (.clk(w377), .nr1(w499), .nr2(w499), .d(w878), .q(w375) );
	dmg_dffr g292 (.clk(w377), .nr1(w499), .nr2(w499), .d(w881), .nq(w881), .q(w814) );
	dmg_dffr g293 (.clk(w164), .nr1(w231), .nr2(w231), .d(w526), .q(w525) );
	dmg_dffr g294 (.clk(w638), .nr1(w386), .nr2(w386), .d(w643), .nq(w643), .q(w644) );
	dmg_dffr g295 (.clk(w643), .nr1(w386), .nr2(w386), .d(w387), .nq(w387), .q(w970) );
	dmg_dffr g296 (.clk(w387), .nr1(w386), .nr2(w386), .d(w579), .nq(w579), .q(w580) );
	dmg_dffr g297 (.clk(w579), .nr1(w386), .nr2(w386), .d(w124), .nq(w124), .q(w125) );
	dmg_dffr g298 (.clk(w124), .nr1(w386), .nr2(w386), .d(w578), .nq(w578), .q(w577) );
	dmg_dffr g299 (.clk(w381), .nr1(w274), .nr2(w274), .d(w275), .nq(w275), .q(w276) );
	dmg_dffr g300 (.clk(w570), .nr1(w274), .nr2(w274), .d(w381), .nq(w381), .q(w382) );
	dmg_dffr g301 (.clk(w568), .nr1(w274), .nr2(w274), .d(w570), .nq(w570), .q(w569) );
	dmg_dffr g302 (.clk(w587), .nr1(w274), .nr2(w274), .d(w568), .nq(w568), .q(w273) );
	dmg_dffr g303 (.clk(w365), .nr1(w148), .nr2(w148), .d(w290), .nq(w290) );
	dmg_dffr g304 (.clk(w364), .nr1(w148), .nr2(w148), .d(w290), .nq(w289), .q(w288) );
	dmg_dffr g305 (.clk(w150), .nr1(w138), .nr2(w138), .d(w149) );
	dmg_dffr g306 (.clk(w44), .nr1(w499), .nr2(w499), .d(w832), .q(w369) );
	dmg_dffr g307 (.clk(w44), .nr1(w499), .nr2(w499), .d(w522), .q(w171) );
	dmg_dffr g308 (.clk(w44), .nr1(w499), .nr2(w499), .d(w498), .nq(w498), .q(w497) );
	dmg_dffr g309 (.clk(w275), .nr1(w274), .nr2(w274), .d(w640), .nq(w640), .q(w639) );
	dmg_dffr g310 (.clk(w800), .nr1(w386), .nr2(w386), .d(w642), .nq(w642), .q(w388) );
	dmg_dffr g311 (.clk(w642), .nr1(w386), .nr2(w386), .d(w385), .nq(w385), .q(w384) );
	dmg_dffr g312 (.clk(w385), .nr1(w386), .nr2(w386), .d(w638), .nq(w638), .q(w334) );
	dmg_dffr g313 (.clk(w319), .nr1(w499), .nr2(w499), .d(w500), .q(w619) );
	dmg_dffr g314 (.clk(w164), .nr1(w231), .nr2(w231), .d(w525), .nq(w243), .q(w242) );
	dmg_dffr g315 (.clk(w290), .nr1(w148), .nr2(w148), .d(w869), .nq(w869) );
	dmg_dffr g316 (.clk(w406), .nr1(w408), .nr2(w408), .d(w407), .nq(w407), .q(w400) );
	dmg_dffr g317 (.clk(w708), .nr1(w408), .nr2(w408), .d(w933), .nq(w933), .q(w706) );
	dmg_dffr g318 (.clk(w975), .nr1(w424), .nr2(w424), .d(w936), .q(w670) );
	dmg_dffr g319 (.clk(w513), .nr1(w408), .nr2(w408), .d(w932), .nq(w932), .q(w404) );
	dmg_dffr g320 (.clk(w513), .nr1(w148), .nr2(w148), .d(w966), .q(w754) );
	dmg_dffr g321 (.clk(w44), .nr1(w499), .nr2(w499), .d(w978), .q(w521) );
	dmg_dffr g322 (.clk(w600), .nr1(w231), .nr2(w231), .d(w242), .q(w230) );
	dmg_dffr g323 (.clk(w377), .nr1(w499), .nr2(w499), .d(w899), .q(w624) );
	dmg_dffr g324 (.clk(w319), .nr1(w148), .nr2(w148), .d(w177), .q(w882) );
	dmg_dffr g325 (.clk(w164), .nr1(w186), .nr2(w186), .d(w876), .q(w185) );
	dmg_dffr g326 (.clk(w600), .nr1(w47), .nr2(w47), .d(w185), .nq(w184) );
	dmg_dffr g327 (.clk(w659), .nr1(w167), .nr2(w167), .d(w875), .q(w179) );
	dmg_dffr g328 (.clk(w319), .nr1(w231), .nr2(w231), .d(w179), .q(w874) );
	dmg_dffr g329 (.clk(w632), .nr1(w231), .nr2(w231), .d(w511), .q(w810) );
	dmg_dffr g330 (.clk(w631), .nr1(w148), .nr2(w148), .d(w628), .q(w168) );
	dmg_dffr g331 (.clk(w632), .nr1(w231), .nr2(w231), .d(w171), .q(w429) );
	dmg_dffr g332 (.clk(w174), .nr1(w424), .nr2(w424), .d(w960), .nq(w740), .q(w739) );
	dmg_dffr g333 (.clk(w173), .nr1(w424), .nr2(w424), .d(w544), .q(w410) );
	dmg_dffr g334 (.clk(w173), .nr1(w424), .nr2(w424), .d(w425), .q(w423) );
	dmg_dffr g335 (.clk(w411), .nr1(w257), .nr2(w257), .d(w493), .nq(w493), .q(w172) );
	dmg_dffr g336 (.clk(w419), .nr1(w257), .nr2(w257), .d(w253), .nq(w253), .q(w252) );
	dmg_dffr g337 (.clk(w253), .nr1(w257), .nr2(w257), .d(w412), .nq(w412), .q(w286) );
	dmg_dffr g338 (.clk(w466), .nr1(w143), .nr2(w143), .d(w465), .nq(w465), .q(w464) );
	dmg_nand g339 (.a(w113), .b(w324), .x(w323) );
	dmg_nand g340 (.a(w326), .b(w113), .x(w762) );
	dmg_nand g341 (.a(w113), .b(w664), .x(w662) );
	dmg_nand g342 (.a(w663), .b(w113), .x(w661) );
	dmg_nand g343 (.a(w113), .b(w331), .x(w329) );
	dmg_nand g344 (.a(w330), .b(w113), .x(w763) );
	dmg_nand g345 (.a(w761), .b(w113), .x(w760) );
	dmg_nand g346 (.a(w113), .b(w317), .x(w316) );
	dmg_nand g347 (.a(w319), .b(w320), .x(w467) );
	dmg_nand g348 (.a(w199), .b(w30), .x(w29) );
	dmg_nand g349 (.a(w947), .b(w30), .x(w977) );
	dmg_nand g350 (.a(w199), .b(w475), .x(w474) );
	dmg_nand g351 (.a(w774), .b(w475), .x(w775) );
	dmg_nand g352 (.a(w28), .b(w438), .x(w938) );
	dmg_nand g353 (.a(w18), .b(w17), .x(w24) );
	dmg_nand g354 (.a(w939), .b(w17), .x(w398) );
	dmg_nand g355 (.a(w27), .b(w438), .x(w399) );
	dmg_nand g356 (.a(w201), .b(w200), .x(w937) );
	dmg_nand g357 (.a(w462), .b(w222), .x(w461) );
	dmg_nand g358 (.a(w113), .b(w328), .x(w759) );
	dmg_nand g359 (.a(w327), .b(w113), .x(w821) );
	dmg_nand g360 (.a(w113), .b(w118), .x(w117) );
	dmg_nand g361 (.a(w315), .b(w113), .x(w758) );
	dmg_nand g362 (.a(w113), .b(w214), .x(w312) );
	dmg_nand g363 (.a(w213), .b(w113), .x(w112) );
	dmg_nand g364 (.a(w142), .b(w46), .x(w581) );
	dmg_nand g365 (.a(w142), .b(w565), .x(w564) );
	dmg_nand g366 (.a(w142), .b(w766), .x(w559) );
	dmg_nand g367 (.a(w588), .b(w142), .x(w141) );
	dmg_nand g368 (.a(w142), .b(w562), .x(w561) );
	dmg_nand g369 (.a(w142), .b(w770), .x(w590) );
	dmg_nand g370 (.a(w142), .b(w858), .x(w591) );
	dmg_nand g371 (.a(w854), .b(w769), .x(w855) );
	dmg_nand g372 (.a(w979), .b(w744), .x(w743) );
	dmg_nand g373 (.a(w669), .b(w21), .x(w782) );
	dmg_nand g374 (.a(w866), .b(w21), .x(w446) );
	dmg_nand g375 (.a(w792), .b(w676), .x(w198) );
	dmg_nand g376 (.a(w199), .b(w676), .x(w675) );
	dmg_nand g377 (.a(w728), .b(w200), .x(w726) );
	dmg_nand g378 (.a(w727), .b(w200), .x(w723) );
	dmg_nand g379 (.a(w793), .b(w200), .x(w731) );
	dmg_nand g380 (.a(w952), .b(w21), .x(w709) );
	dmg_nand g381 (.a(w716), .b(w676), .x(w677) );
	dmg_nand g382 (.a(w717), .b(w17), .x(w718) );
	dmg_nand g383 (.a(w527), .b(w17), .x(w931) );
	dmg_nand g384 (.a(w953), .b(w475), .x(w476) );
	dmg_nand g385 (.a(w308), .b(w307), .x(w955) );
	dmg_nand g386 (.a(w691), .b(w307), .x(w690) );
	dmg_nand g387 (.a(w33), .b(w307), .x(w692) );
	dmg_nand g388 (.a(w872), .b(w307), .x(w954) );
	dmg_nand g389 (.a(w306), .b(w30), .x(w871) );
	dmg_nand g390 (.a(w35), .b(w30), .x(w870) );
	dmg_nand g391 (.a(w527), .b(w307), .x(w301) );
	dmg_nand g392 (.a(w527), .b(w30), .x(w299) );
	dmg_nand g393 (.a(w527), .b(w188), .x(w187) );
	dmg_nand g394 (.a(w868), .b(w205), .x(w206) );
	dmg_nand g395 (.a(w227), .b(w229), .x(w599) );
	dmg_nand g396 (.a(w882), .b(w656), .x(w501) );
	dmg_nand g397 (.a(w688), .b(w30), .x(w689) );
	dmg_nand g398 (.a(w686), .b(w188), .x(w189) );
	dmg_nand g399 (.a(w841), .b(w195), .x(w685) );
	dmg_nand g400 (.a(w839), .b(w21), .x(w934) );
	dmg_nand g401 (.a(w713), .b(w676), .x(w715) );
	dmg_nand g402 (.a(w956), .b(w676), .x(w959) );
	dmg_nand g403 (.a(w833), .b(w200), .x(w681) );
	dmg_nand g404 (.a(w527), .b(w200), .x(w680) );
	dmg_nand g405 (.a(w527), .b(w676), .x(w683) );
	dmg_nand g406 (.a(w527), .b(w21), .x(w928) );
	dmg_nand g407 (.a(w714), .b(w676), .x(w840) );
	dmg_nand g408 (.a(w304), .b(w195), .x(w929) );
	dmg_nand g409 (.a(w830), .b(w195), .x(w845) );
	dmg_nand g410 (.a(w842), .b(w30), .x(w843) );
	dmg_nand g411 (.a(w527), .b(w195), .x(w303) );
	dmg_nand g412 (.a(w81), .b(w82), .x(w961) );
	dmg_nand g413 (.a(w210), .b(w145), .x(w383) );
	dmg_nand g414 (.a(w603), .b(w30), .x(w478) );
	dmg_nand g415 (.a(w32), .b(w195), .x(w844) );
	dmg_nand g416 (.a(w305), .b(w195), .x(w192) );
	dmg_nand g417 (.a(w488), .b(w676), .x(w720) );
	dmg_nand g418 (.a(w199), .b(w200), .x(w730) );
	dmg_nand g419 (.a(w199), .b(w21), .x(w710) );
	dmg_nand g420 (.a(w867), .b(w188), .x(w671) );
	dmg_nand g421 (.a(w600), .b(w599), .x(w822) );
	dmg_nand g422 (.a(w917), .b(w142), .x(w912) );
	dmg_nand g423 (.a(w913), .b(w142), .x(w908) );
	dmg_nand g424 (.a(w556), .b(w142), .x(w768) );
	dmg_nand g425 (.a(w142), .b(w767), .x(w910) );
	dmg_nand g426 (.a(w860), .b(w142), .x(w911) );
	dmg_nand g427 (.a(w967), .b(w142), .x(w918) );
	dmg_nand g428 (.a(w969), .b(w142), .x(w968) );
	dmg_nand g429 (.a(w45), .b(w142), .x(w557) );
	dmg_nand g430 (.a(w632), .b(w507), .x(w506) );
	dmg_nand g431 (.a(w199), .b(w188), .x(w945) );
	dmg_nand g432 (.a(w447), .b(w188), .x(w942) );
	dmg_nand g433 (.a(w199), .b(w17), .x(w674) );
	dmg_nand g434 (.a(w528), .b(w17), .x(w790) );
	dmg_nand g435 (.a(w444), .b(w17), .x(w724) );
	dmg_nand g436 (.a(w16), .b(w17), .x(w725) );
	dmg_nand g437 (.a(w202), .b(w200), .x(w805) );
	dmg_nand g438 (.a(w487), .b(w21), .x(w788) );
	dmg_nand g439 (.a(w20), .b(w21), .x(w785) );
	dmg_nand g440 (.a(w437), .b(w188), .x(w941) );
	dmg_nand g441 (.a(w19), .b(w188), .x(w15) );
	dmg_nand g442 (.a(w199), .b(w195), .x(w196) );
	dmg_nand g443 (.a(w925), .b(w113), .x(w114) );
	dmg_nand g444 (.a(w113), .b(w216), .x(w215) );
	dmg_latch_comp g445 (.n_ena(w219), .d(w218), .ena(w119), .q(w324) );
	dmg_latch_comp g446 (.n_ena(w219), .d(w332), .ena(w119), .q(w331) );
	dmg_latch_comp g447 (.n_ena(w219), .d(w553), .ena(w119), .q(w328) );
	dmg_latch_comp g448 (.n_ena(w219), .d(w554), .ena(w119), .q(w118) );
	dmg_latch_comp g449 (.n_ena(w219), .d(w120), .ena(w119), .q(w214) );
	dmg_latch_comp g450 (.n_ena(w449), .d(w310), .ena(w34), .q(w35) );
	dmg_latch_comp g451 (.n_ena(w449), .d(w450), .ena(w34), .q(w33) );
	dmg_latch_comp g452 (.n_ena(w449), .d(w448), .ena(w34), .q(w728) );
	dmg_latch_comp g453 (.n_ena(w451), .d(w886), .ena(w309), .q(w447) );
	dmg_latch_comp g454 (.n_ena(w449), .d(w771), .ena(w34), .q(w669) );
	dmg_latch_comp g455 (.n_ena(w451), .d(w489), .ena(w309), .q(w488) );
	dmg_latch_comp g456 (.n_ena(w449), .d(w489), .ena(w34), .q(w716) );
	dmg_latch_comp g457 (.n_ena(w451), .d(w450), .ena(w309), .q(w308) );
	dmg_latch_comp g458 (.n_ena(w449), .d(w873), .ena(w34), .q(w32) );
	dmg_latch_comp g459 (.n_ena(w451), .d(w873), .ena(w309), .q(w305) );
	dmg_latch_comp g460 (.n_ena(w451), .d(w310), .ena(w309), .q(w603) );
	dmg_latch_comp g461 (.n_ena(w451), .d(w448), .ena(w309), .q(w202) );
	dmg_latch_comp g462 (.n_ena(w449), .d(w886), .ena(w34), .q(w19) );
	dmg_latch_comp g463 (.n_ena(w451), .d(w771), .ena(w309), .q(w20) );
	dmg_latch_comp g464 (.n_ena(w451), .d(w459), .ena(w309), .q(w18) );
	dmg_latch_comp g465 (.n_ena(w449), .d(w459), .ena(w34), .q(w16) );
	dmg_latch_comp g466 (.n_ena(w219), .d(w121), .ena(w119), .q(w317) );
	dmg_latch_comp g467 (.n_ena(w219), .d(w217), .ena(w119), .q(w216) );
	dmg_latch_comp g468 (.n_ena(w219), .d(w311), .ena(w119), .q(w664) );
	dmg_not2 g469 (.a(w325), .x(w212) );
	dmg_not2 g470 (.a(w665), .x(w314) );
	dmg_not2 g471 (.a(w314), .x(w313) );
	dmg_not2 g472 (.a(w143), .x(w142) );
	dmg_not2 g473 (.a(w143), .x(w113) );
	dmg_not2 g474 (.a(w389), .x(w390) );
	dmg_not2 g475 (.a(w518), .x(w471) );
	dmg_not2 g476 (.a(w515), .x(w514) );
	dmg_not2 g477 (.a(w801), .x(w802) );
	dmg_not2 g478 (.a(w50), .x(w51) );
	dmg_not2 g479 (.a(w895), .x(w472) );
	dmg_not2 g480 (.a(w155), .x(w156) );
	dmg_not2 g481 (.a(w278), .x(w279) );
	dmg_not2 g482 (.a(w61), .x(w62) );
	dmg_not2 g483 (.a(w3), .x(w4) );
	dmg_not2 g484 (.a(w529), .x(w530) );
	dmg_not2 g485 (.a(w586), .x(w585) );
	dmg_not2 g486 (.a(w797), .x(w796) );
	dmg_not2 g487 (.a(w163), .x(w877) );
	dmg_nand g488 (.a(w142), .x(w914), .b(w596) );
	dmg_not2 g489 (.a(w597), .x(w123) );
	dmg_not2 g490 (.a(w516), .x(w576) );
	dmg_not2 g491 (.a(w572), .x(w268) );
	dmg_not2 g492 (.a(w649), .x(w650) );
	dmg_not2 g493 (.a(w137), .x(w250) );
	dmg_not2 g494 (.a(w292), .x(w293) );
	dmg_not2 g495 (.a(w137), .x(w247) );
	dmg_not2 g496 (.a(w848), .x(w847) );
	dmg_not2 g497 (.a(w961), .x(w148) );
	dmg_not2 g498 (.a(w288), .x(w287) );
	dmg_not2 g499 (.a(w290), .x(w496) );
	dmg_not2 g500 (.a(w75), .x(w74) );
	dmg_not2 g501 (.a(w243), .x(w244) );
	dmg_not2 g502 (.a(w920), .x(w73) );
	dmg_not2 g503 (.a(w849), .x(w850) );
	dmg_not2 g504 (.a(w263), .x(w262) );
	dmg_not2 g505 (.a(w269), .x(w270) );
	dmg_not2 g506 (.a(w136), .x(w137) );
	dmg_not2 g507 (.a(w238), .x(w237) );
	dmg_not2 g508 (.a(w571), .x(w641) );
	dmg_not2 g509 (.a(w161), .x(w160) );
	dmg_not2 g510 (.a(w798), .x(w537) );
	dmg_not2 g511 (.a(w235), .x(w234) );
	dmg_not2 g512 (.a(w926), .x(w294) );
	dmg_not2 g513 (.a(w781), .x(w687) );
	dmg_not2 g514 (.a(w855), .x(w824) );
	dmg_not2 g515 (.a(w501), .x(w905) );
	dmg_not2 g516 (.a(w146), .x(w145) );
	dmg_not2 g517 (.a(w865), .x(w950) );
	dmg_not2 g518 (.a(w64), .x(w63) );
	dmg_not2 g519 (.a(w583), .x(w584) );
	dmg_not2 g520 (.a(w808), .x(w898) );
	dmg_notif0 g521 (.n_ena(w95), .a(w434), .x(w341) );
	dmg_notif0 g522 (.n_ena(w95), .a(w863), .x(w13) );
	dmg_notif0 g523 (.n_ena(w95), .a(w96), .x(w91) );
	dmg_notif0 g524 (.n_ena(w95), .a(w803), .x(w79) );
	dmg_notif0 g525 (.n_ena(w95), .a(w896), .x(w249) );
	dmg_notif0 g526 (.n_ena(w95), .a(w100), .x(w52) );
	dmg_notif0 g527 (.n_ena(w95), .a(w94), .x(w68) );
	dmg_notif0 g528 (.n_ena(w95), .a(w890), .x(w12) );
	dmg_notif0 g529 (.n_ena(w372), .a(w519), .x(w13) );
	dmg_notif0 g530 (.n_ena(w372), .a(w892), .x(w52) );
	dmg_notif0 g531 (.n_ena(w260), .a(w259), .x(w91) );
	dmg_notif0 g532 (.n_ena(w158), .a(w157), .x(w52) );
	dmg_notif0 g533 (.n_ena(w453), .a(w101), .x(w52) );
	dmg_notif0 g534 (.n_ena(w453), .a(w734), .x(w68) );
	dmg_notif0 g535 (.n_ena(w453), .a(w735), .x(w79) );
	dmg_notif0 g536 (.n_ena(w453), .a(w492), .x(w341) );
	dmg_notif0 g537 (.n_ena(w453), .a(w484), .x(w249) );
	dmg_notif0 g538 (.n_ena(w237), .a(w593), .x(w48) );
	dmg_notif0 g539 (.n_ena(w237), .a(w594), .x(w566) );
	dmg_notif0 g540 (.n_ena(w237), .a(w333), .x(w126) );
	dmg_notif0 g541 (.n_ena(w237), .a(w595), .x(w60) );
	dmg_notif0 g542 (.n_ena(w237), .a(w555), .x(w65) );
	dmg_notif0 g543 (.n_ena(w67), .a(w752), .x(w91) );
	dmg_notif0 g544 (.n_ena(w67), .a(w751), .x(w13) );
	dmg_notif0 g545 (.n_ena(w67), .a(w606), .x(w52) );
	dmg_notif0 g546 (.n_ena(w67), .a(w605), .x(w68) );
	dmg_notif0 g547 (.n_ena(w453), .a(w107), .x(w13) );
	dmg_notif0 g548 (.n_ena(w453), .a(w452), .x(w91) );
	dmg_notif0 g549 (.n_ena(w383), .a(w384), .x(w154) );
	dmg_notif0 g550 (.n_ena(w335), .a(w388), .x(w131) );
	dmg_notif0 g551 (.n_ena(w335), .a(w334), .x(w277) );
	dmg_notif0 g552 (.n_ena(w576), .a(w639), .x(w517) );
	dmg_notif0 g553 (.n_ena(w57), .a(w86), .x(w13) );
	dmg_notif0 g554 (.n_ena(w57), .a(w53), .x(w52) );
	dmg_notif0 g555 (.n_ena(w57), .a(w56), .x(w91) );
	dmg_notif0 g556 (.n_ena(w284), .a(w337), .x(w249) );
	dmg_notif0 g557 (.n_ena(w284), .a(w78), .x(w79) );
	dmg_notif0 g558 (.n_ena(w284), .a(w338), .x(w52) );
	dmg_notif0 g559 (.n_ena(w284), .a(w360), .x(w341) );
	dmg_notif0 g560 (.n_ena(w284), .a(w285), .x(w12) );
	dmg_notif0 g561 (.n_ena(w343), .a(w344), .x(w13) );
	dmg_notif0 g562 (.n_ena(w343), .a(w958), .x(w91) );
	dmg_notif0 g563 (.n_ena(w343), .a(w359), .x(w52) );
	dmg_notif0 g564 (.n_ena(w343), .a(w350), .x(w79) );
	dmg_notif0 g565 (.n_ena(w343), .a(w342), .x(w341) );
	dmg_notif0 g566 (.n_ena(w343), .a(w831), .x(w249) );
	dmg_notif0 g567 (.n_ena(w343), .a(w836), .x(w68) );
	dmg_notif0 g568 (.n_ena(w343), .a(w835), .x(w12) );
	dmg_notif0 g569 (.n_ena(w57), .a(w980), .x(w12) );
	dmg_notif0 g570 (.n_ena(w57), .a(w80), .x(w79) );
	dmg_notif0 g571 (.n_ena(w237), .a(w133), .x(w49) );
	dmg_notif0 g572 (.n_ena(w237), .a(w132), .x(w154) );
	dmg_notif0 g573 (.n_ena(w237), .a(w574), .x(w517) );
	dmg_notif0 g574 (.n_ena(w237), .a(w134), .x(w135) );
	dmg_notif0 g575 (.n_ena(w237), .a(w127), .x(w271) );
	dmg_notif0 g576 (.n_ena(w335), .a(w223), .x(w272) );
	dmg_notif0 g577 (.n_ena(w237), .a(w919), .x(w272) );
	dmg_notif0 g578 (.n_ena(w237), .a(w130), .x(w131) );
	dmg_notif0 g579 (.n_ena(w576), .a(w273), .x(w272) );
	dmg_notif0 g580 (.n_ena(w237), .a(w129), .x(w277) );
	dmg_notif0 g581 (.n_ena(w576), .a(w569), .x(w131) );
	dmg_notif0 g582 (.n_ena(w576), .a(w382), .x(w154) );
	dmg_notif0 g583 (.n_ena(w576), .a(w276), .x(w277) );
	dmg_notif0 g584 (.n_ena(w576), .a(w577), .x(w566) );
	dmg_notif0 g585 (.n_ena(w576), .a(w125), .x(w126) );
	dmg_notif0 g586 (.n_ena(w576), .a(w580), .x(w135) );
	dmg_notif0 g587 (.n_ena(w576), .a(w970), .x(w271) );
	dmg_notif0 g588 (.n_ena(w576), .a(w644), .x(w49) );
	dmg_notif0 g589 (.n_ena(w576), .a(w47), .x(w48) );
	dmg_notif0 g590 (.n_ena(w576), .a(w645), .x(w60) );
	dmg_notif0 g591 (.n_ena(w576), .a(w47), .x(w65) );
	dmg_notif0 g592 (.n_ena(w57), .a(w540), .x(w249) );
	dmg_notif0 g593 (.n_ena(w57), .a(w87), .x(w68) );
	dmg_notif0 g594 (.n_ena(w57), .a(w880), .x(w341) );
	dmg_notif0 g595 (.n_ena(w67), .a(w66), .x(w12) );
	dmg_notif0 g596 (.n_ena(w260), .a(w974), .x(w68) );
	dmg_notif0 g597 (.n_ena(w260), .a(w973), .x(w13) );
	dmg_notif0 g598 (.n_ena(w67), .a(w291), .x(w249) );
	dmg_notif0 g599 (.n_ena(w67), .a(w753), .x(w341) );
	dmg_notif0 g600 (.n_ena(w479), .a(w857), .x(w341) );
	dmg_notif0 g601 (.n_ena(w158), .a(w428), .x(w12) );
	dmg_notif0 g602 (.n_ena(w67), .a(w430), .x(w79) );
	dmg_notif0 g603 (.n_ena(w158), .a(w90), .x(w91) );
	dmg_notif0 g604 (.n_ena(w158), .a(w547), .x(w249) );
	dmg_notif0 g605 (.n_ena(w158), .a(w512), .x(w13) );
	dmg_notif0 g606 (.n_ena(w158), .a(w433), .x(w341) );
	dmg_notif0 g607 (.n_ena(w479), .a(w480), .x(w68) );
	dmg_notif0 g608 (.n_ena(w479), .a(w548), .x(w249) );
	dmg_notif0 g609 (.n_ena(w479), .a(w483), .x(w52) );
	dmg_notif0 g610 (.n_ena(w453), .a(w454), .x(w12) );
	dmg_notif0 g611 (.n_ena(w158), .a(w494), .x(w68) );
	dmg_notif0 g612 (.n_ena(w158), .a(w283), .x(w79) );
	dmg_notif0 g613 (.n_ena(w372), .a(w371), .x(w91) );
	dmg_notif0 g614 (.n_ena(w372), .a(w891), .x(w341) );
	dmg_notif0 g615 (.n_ena(w372), .a(w812), .x(w79) );
	dmg_notif0 g616 (.n_ena(w372), .a(w820), .x(w68) );
	dmg_notif0 g617 (.n_ena(w372), .a(w373), .x(w249) );
	dmg_notif0 g618 (.n_ena(w372), .a(w646), .x(w12) );
	dmg_latchnq_comp g619 (.n_ena(w93), .d(w79), .ena(w92), .q(w804), .nq(w803) );
	dmg_latchnq_comp g620 (.n_ena(w93), .d(w341), .ena(w92), .q(w435), .nq(w434) );
	dmg_latchnq_comp g621 (.n_ena(w93), .d(w249), .ena(w92), .q(w391), .nq(w896) );
	dmg_latchnq_comp g622 (.n_ena(w93), .d(w52), .ena(w92), .q(w99), .nq(w100) );
	dmg_latchnq_comp g623 (.n_ena(w93), .d(w68), .ena(w92), .q(w806), .nq(w94) );
	dmg_latchnq_comp g624 (.n_ena(w93), .d(w12), .ena(w92), .q(w889), .nq(w890) );
	dmg_latchnq_comp g625 (.n_ena(w108), .d(w12), .ena(w733), .q(w455), .nq(w454) );
	dmg_latchnq_comp g626 (.n_ena(w69), .d(w12), .ena(w70), .q(w834), .nq(w835) );
	dmg_latchnq_comp g627 (.n_ena(w69), .d(w68), .ena(w70), .q(w837), .nq(w836) );
	dmg_latchnq_comp g628 (.n_ena(w69), .d(w249), .ena(w70), .q(w838), .nq(w831) );
	dmg_latchnq_comp g629 (.n_ena(w69), .d(w341), .ena(w70), .q(w349), .nq(w342) );
	dmg_latchnq_comp g630 (.n_ena(w69), .d(w79), .ena(w70), .q(w351), .nq(w350) );
	dmg_latchnq_comp g631 (.n_ena(w69), .d(w52), .ena(w70), .q(w358), .nq(w359) );
	dmg_latchnq_comp g632 (.n_ena(w69), .d(w91), .ena(w70), .q(w957), .nq(w958) );
	dmg_latchnq_comp g633 (.n_ena(w69), .d(w13), .ena(w70), .q(w345), .nq(w344) );
	dmg_latchr_comp g634 (.n_ena(w88), .d(w79), .ena(w818), .nres(w250), .q(w811), .nq(w812) );
	dmg_latchr_comp g635 (.n_ena(w88), .d(w12), .ena(w818), .nres(w250), .q(w647), .nq(w646) );
	dmg_latchr_comp g636 (.n_ena(w88), .d(w91), .ena(w818), .nres(w250), .q(w370), .nq(w371) );
	dmg_latchr_comp g637 (.n_ena(w295), .d(w79), .ena(w413), .nres(w250), .q(w282), .nq(w283) );
	dmg_latchr_comp g638 (.n_ena(w295), .d(w12), .ena(w413), .nres(w250), .q(w416), .nq(w428) );
	dmg_latchr_comp g639 (.n_ena(w295), .d(w91), .ena(w413), .nres(w250), .q(w89), .nq(w90) );
	dmg_latchr_comp g640 (.n_ena(w295), .d(w68), .ena(w413), .nres(w250), .q(w495), .nq(w494) );
	dmg_latchr_comp g641 (.n_ena(w295), .d(w249), .ena(w413), .nres(w250), .q(w546), .nq(w547) );
	dmg_latchr_comp g642 (.n_ena(w295), .d(w341), .ena(w413), .nres(w250), .q(w545), .nq(w433) );
	dmg_latchr_comp g643 (.n_ena(w295), .d(w13), .ena(w413), .nres(w250), .q(w251), .nq(w512) );
	dmg_latchr_comp g644 (.n_ena(w613), .d(w341), .ena(w612), .nres(w247), .q(w779), .nq(w857) );
	dmg_latchr_comp g645 (.n_ena(w613), .d(w68), .ena(w612), .nres(w247), .q(w481), .nq(w480) );
	dmg_latchr_comp g646 (.n_ena(w613), .d(w52), .ena(w612), .nres(w247), .q(w482), .nq(w483) );
	dmg_latchr_comp g647 (.n_ena(w613), .d(w249), .ena(w612), .nres(w247), .q(w549), .nq(w548) );
	dmg_latchr_comp g648 (.n_ena(w71), .d(w79), .ena(w248), .nres(w247), .q(w611), .nq(w430) );
	dmg_latchr_comp g649 (.n_ena(w85), .d(w249), .ena(w539), .nres(w138), .q(w645), .nq(w540) );
	dmg_latchr_comp g650 (.n_ena(w85), .d(w68), .ena(w539), .nres(w138), .q(w208), .nq(w87) );
	dmg_latchr_comp g651 (.n_ena(w85), .d(w341), .ena(w539), .nres(w138), .q(w542), .nq(w880) );
	dmg_latchr_comp g652 (.n_ena(w83), .d(w79), .ena(w84), .nres(w82), .q(w149) );
	dmg_latchr_comp g653 (.n_ena(w85), .d(w91), .ena(w539), .nres(w138), .q(w55), .nq(w56) );
	dmg_latchr_comp g654 (.n_ena(w85), .d(w52), .ena(w539), .nres(w138), .q(w54), .nq(w53) );
	dmg_latchr_comp g655 (.n_ena(w85), .d(w12), .ena(w539), .nres(w138), .q(w829), .nq(w980) );
	dmg_latchr_comp g656 (.n_ena(w85), .d(w79), .ena(w539), .nres(w138), .q(w81), .nq(w80) );
	dmg_latchr_comp g657 (.n_ena(w85), .d(w13), .ena(w539), .nres(w138), .q(w139), .nq(w86) );
	dmg_latchr_comp g658 (.n_ena(w71), .d(w12), .ena(w248), .nres(w247), .q(w856), .nq(w66) );
	dmg_latchr_comp g659 (.n_ena(w71), .d(w341), .ena(w248), .nres(w247), .q(w879), .nq(w753) );
	dmg_latchr_comp g660 (.n_ena(w71), .d(w249), .ena(w248), .nres(w247), .q(w608), .nq(w291) );
	dmg_latchr_comp g661 (.n_ena(w71), .d(w68), .ena(w248), .nres(w247), .q(w604), .nq(w605) );
	dmg_latchr_comp g662 (.n_ena(w71), .d(w52), .ena(w248), .nres(w247), .q(w607), .nq(w606) );
	dmg_latchr_comp g663 (.n_ena(w71), .d(w13), .ena(w248), .nres(w247), .q(w750), .nq(w751) );
	dmg_latchr_comp g664 (.n_ena(w71), .d(w91), .ena(w248), .nres(w247), .q(w246), .nq(w752) );
	dmg_latchr_comp g665 (.n_ena(w295), .d(w52), .ena(w413), .nres(w250), .q(w254), .nq(w157) );
	dmg_latchr_comp g666 (.n_ena(w88), .d(w52), .ena(w818), .nres(w250), .q(w893), .nq(w892) );
	dmg_latchr_comp g667 (.n_ena(w88), .d(w341), .ena(w818), .nres(w250), .q(w964), .nq(w891) );
	dmg_latchr_comp g668 (.n_ena(w88), .d(w13), .ena(w818), .nres(w250), .q(w520), .nq(w519) );
	dmg_latchr_comp g669 (.n_ena(w88), .d(w249), .ena(w818), .nres(w250), .q(w374), .nq(w373) );
	dmg_latchr_comp g670 (.n_ena(w88), .d(w68), .ena(w818), .nres(w250), .q(w813), .nq(w820) );
	dmg_latchnq_comp g671 (.n_ena(w93), .d(w13), .ena(w92), .q(w864), .nq(w863) );
	dmg_latchnq_comp g672 (.n_ena(w93), .d(w91), .ena(w92), .q(w97), .nq(w96) );
	dmg_latchnq_comp g673 (.n_ena(w108), .d(w52), .ena(w733), .q(w102), .nq(w101) );
	dmg_latchnq_comp g674 (.n_ena(w108), .d(w68), .ena(w733), .q(w737), .nq(w734) );
	dmg_latchnq_comp g675 (.n_ena(w108), .d(w79), .ena(w733), .q(w736), .nq(w735) );
	dmg_latchnq_comp g676 (.n_ena(w108), .d(w341), .ena(w733), .q(w491), .nq(w492) );
	dmg_latchnq_comp g677 (.n_ena(w108), .d(w249), .ena(w733), .q(w485), .nq(w484) );
	dmg_latchnq_comp g678 (.n_ena(w108), .d(w91), .ena(w733), .q(w490), .nq(w452) );
	dmg_latchnq_comp g679 (.n_ena(w108), .d(w13), .ena(w733), .q(w106), .nq(w107) );
	dmg_nand g680 (.a(w943), .b(w188), .x(w787) );
	dmg_nand g681 (.a(w951), .b(w195), .x(w777) );
	dmg_and g682 (.a(w318), .b(w231), .x(w660) );
	dmg_and g683 (.a(w461), .b(w212), .x(w210) );
	dmg_and g684 (.a(w462), .b(w463), .x(w666) );
	dmg_and g685 (.a(w59), .b(w877), .x(w862) );
	dmg_and g686 (.a(w152), .b(w877), .x(w807) );
	dmg_and g687 (.a(w460), .b(w212), .x(w211) );
	dmg_and g688 (.a(w147), .b(w634), .x(w633) );
	dmg_and g689 (.a(w809), .b(w810), .x(w7) );
	dmg_and g690 (.a(w242), .b(w204), .x(w203) );
	dmg_and g691 (.a(w526), .b(w204), .x(w693) );
	dmg_and g692 (.a(w59), .b(w234), .x(w233) );
	dmg_and g693 (.a(w207), .b(w687), .x(w780) );
	dmg_and g694 (.a(w668), .b(w298), .x(w439) );
	dmg_and g695 (.a(w297), .b(w298), .x(w440) );
	dmg_and g696 (.a(w152), .b(w234), .x(w601) );
	dmg_and g697 (.a(w376), .b(w375), .x(w900) );
	dmg_and g698 (.a(w500), .b(w207), .x(w655) );
	dmg_and g699 (.a(w524), .b(w44), .x(w903) );
	dmg_and g700 (.a(w756), .b(w139), .x(w668) );
	dmg_and g701 (.a(w184), .b(w185), .x(w534) );
	dmg_and g702 (.a(w206), .b(w123), .x(w582) );
	dmg_and g703 (.a(w211), .b(w145), .x(w516) );
	dmg_and g704 (.a(w144), .b(w145), .x(w587) );
	dmg_and g705 (.a(w153), .b(w123), .x(w122) );
	dmg_and g706 (.a(w59), .b(w537), .x(w921) );
	dmg_and g707 (.a(w621), .b(w622), .x(w500) );
	dmg_and g708 (.a(w497), .b(w171), .x(w523) );
	dmg_and g709 (.a(w206), .b(w226), .x(w225) );
	dmg_and g710 (.a(w152), .b(w537), .x(w538) );
	dmg_and g711 (.a(w59), .b(w262), .x(w261) );
	dmg_and g712 (.a(w294), .b(w59), .x(w58) );
	dmg_and g713 (.a(w152), .b(w160), .x(w296) );
	dmg_and g714 (.a(w59), .b(w160), .x(w159) );
	dmg_and g715 (.a(w152), .b(w650), .x(w109) );
	dmg_and g716 (.a(w59), .b(w650), .x(w651) );
	dmg_and g717 (.a(w294), .b(w152), .x(w84) );
	dmg_and g718 (.a(w59), .b(w73), .x(w927) );
	dmg_and g719 (.a(w852), .b(w369), .x(w617) );
	dmg_and g720 (.a(w497), .b(w521), .x(w852) );
	dmg_and g721 (.a(w814), .b(w551), .x(w376) );
	dmg_and g722 (.a(w226), .b(w240), .x(w340) );
	dmg_and g723 (.a(w824), .b(w152), .x(w151) );
	dmg_and g724 (.a(w152), .b(w73), .x(w72) );
	dmg_and g725 (.a(w281), .b(w77), .x(w960) );
	dmg_and g726 (.a(w59), .b(w847), .x(w962) );
	dmg_and g727 (.a(w152), .b(w847), .x(w846) );
	dmg_and g728 (.a(w829), .b(w43), .x(w442) );
	dmg_and g729 (.a(w829), .b(w42), .x(w699) );
	dmg_xnor g730 (.b(w813), .a(w814), .x(w635) );
	dmg_xnor g731 (.b(w374), .a(w375), .x(w817) );
	dmg_xnor g732 (.b(w964), .a(w815), .x(w816) );
	dmg_xnor g733 (.b(w893), .a(w171), .x(w170) );
	dmg_xnor g734 (.b(w255), .a(w254), .x(w414) );
	dmg_xnor g735 (.b(w77), .a(w282), .x(w427) );
	dmg_xnor g736 (.b(w281), .a(w495), .x(w543) );
	dmg_xnor g737 (.b(w252), .a(w251), .x(w432) );
	dmg_xnor g738 (.b(w883), .a(w828), .x(w827) );
	dmg_xnor g739 (.b(w508), .a(w11), .x(w10) );
	dmg_xnor g740 (.b(w884), .a(w825), .x(w826) );
	dmg_xnor g741 (.b(w811), .a(w624), .x(w625) );
	dmg_xnor g742 (.b(w647), .a(w521), .x(w948) );
	dmg_xnor g743 (.b(w520), .a(w497), .x(w894) );
	dmg_xnor g744 (.b(w370), .a(w369), .x(w169) );
	dmg_xnor g745 (.b(w286), .a(w416), .x(w431) );
	dmg_xnor g746 (.b(w245), .a(w89), .x(w415) );
	dmg_xnor g747 (.b(w172), .a(w546), .x(w748) );
	dmg_xnor g748 (.b(w361), .a(w545), .x(w747) );
	dmg_nand3 g749 (.a(w463), .b(w464), .c(w222), .x(w221) );
	dmg_nand3 g750 (.a(w861), .b(w143), .c(w468), .x(w320) );
	dmg_nand3 g751 (.a(w229), .b(w230), .c(w242), .x(w241) );
	dmg_nand3 g752 (.a(w883), .b(w884), .c(w508), .x(w507) );
	dmg_nand3 g753 (.a(w128), .b(w127), .c(w573), .x(w572) );
	dmg_nand3 g754 (.a(w542), .b(w541), .c(w148), .x(w336) );
	dmg_not g755 (.a(w488), .x(w714) );
	dmg_and3 g756 (.a(w789), .b(w394), .c(w393), .x(w1) );
	dmg_and3 g757 (.a(w396), .b(w397), .c(w393), .x(w98) );
	dmg_and3 g758 (.a(w395), .b(w397), .c(w393), .x(w26) );
	dmg_and3 g759 (.a(w395), .b(w394), .c(w393), .x(w392) );
	dmg_and3 g760 (.a(w111), .b(w458), .c(w104), .x(w456) );
	dmg_and3 g761 (.a(w110), .b(w457), .c(w104), .x(w103) );
	dmg_and3 g762 (.a(w111), .b(w457), .c(w104), .x(w486) );
	dmg_and3 g763 (.a(w110), .b(w458), .c(w104), .x(w105) );
	dmg_and3 g764 (.a(w502), .b(w503), .c(w915), .x(w904) );
	dmg_and3 g765 (.a(w354), .b(w353), .c(w347), .x(w352) );
	dmg_and3 g766 (.a(w356), .b(w353), .c(w347), .x(w357) );
	dmg_and3 g767 (.a(w354), .b(w355), .c(w347), .x(w348) );
	dmg_and3 g768 (.a(w356), .b(w355), .c(w347), .x(w346) );
	dmg_nor g769 (.a(w699), .b(w442), .x(w441) );
	dmg_nor g770 (.a(w419), .b(w409), .x(w408) );
	dmg_nor g771 (.a(w410), .b(w409), .x(w257) );
	dmg_nor g772 (.a(w533), .b(w532), .x(w653) );
	dmg_nor g773 (.a(w633), .b(w177), .x(w178) );
	dmg_nor g774 (.a(w507), .b(w628), .x(w629) );
	dmg_nor g775 (.a(w667), .b(w898), .x(w167) );
	dmg_nor g776 (.a(w575), .b(w231), .x(w238) );
	dmg_nor g777 (.a(w562), .b(w208), .x(w209) );
	dmg_nor g778 (.a(w916), .b(w907), .x(w906) );
	dmg_nor g779 (.a(w851), .b(w648), .x(w499) );
	dmg_nor g780 (.a(w289), .b(w290), .x(w363) );
	dmg_nor g781 (.a(w368), .b(w231), .x(w239) );
	dmg_nor g782 (.a(w231), .b(w175), .x(w232) );
	dmg_nor g783 (.a(w526), .b(w242), .x(w652) );
	dmg_nand7 g784 (.a(w704), .b(w707), .c(w702), .d(w935), .e(w400), .f(w794), .g(w404), .x(w403) );
	dmg_nand7 g785 (.a(w704), .b(w703), .c(w702), .d(w401), .e(w400), .f(w405), .g(w404), .x(w701) );
	dmg_nand7 g786 (.a(w711), .b(w703), .c(w706), .d(w401), .e(w705), .f(w405), .g(w404), .x(w402) );
	dmg_nand7 g787 (.a(w704), .b(w703), .c(w702), .d(w401), .e(w705), .f(w794), .g(w795), .x(w700) );
	dmg_nand5 g788 (.a(w268), .b(w267), .c(w265), .d(w264), .e(w236), .x(w571) );
	dmg_nand5 g789 (.a(w268), .b(w267), .c(w265), .d(w799), .e(w236), .x(w269) );
	dmg_nand5 g790 (.a(w268), .b(w267), .c(w567), .d(w799), .e(w162), .x(w848) );
	dmg_nand5 g791 (.a(w268), .b(w267), .c(w567), .d(w264), .e(w236), .x(w263) );
	dmg_nand5 g792 (.a(w268), .b(w266), .c(w265), .d(w799), .e(w162), .x(w798) );
	dmg_nand5 g793 (.a(w268), .b(w267), .c(w265), .d(w799), .e(w162), .x(w161) );
	dmg_nand5 g794 (.a(w268), .b(w267), .c(w567), .d(w799), .e(w236), .x(w926) );
	dmg_nand5 g795 (.a(w268), .b(w266), .c(w567), .d(w799), .e(w236), .x(w235) );
	dmg_nand5 g796 (.a(w268), .b(w266), .c(w265), .d(w799), .e(w236), .x(w849) );
	dmg_nand5 g797 (.a(w268), .b(w266), .c(w567), .d(w264), .e(w236), .x(w920) );
	dmg_nand5 g798 (.a(w268), .b(w266), .c(w265), .d(w264), .e(w236), .x(w649) );
	dmg_nand5 g799 (.a(w497), .b(w521), .c(w369), .d(w551), .e(w624), .x(w623) );
	dmg_nand5 g800 (.a(w268), .b(w266), .c(w567), .d(w799), .e(w162), .x(w163) );
	dmg_nand5 g801 (.a(w636), .b(w635), .c(w816), .d(w817), .e(w625), .x(w626) );
	dmg_nand5 g802 (.a(w749), .b(w432), .c(w431), .d(w415), .e(w414), .x(w965) );
	dmg_nand5 g803 (.a(w542), .b(w543), .c(w747), .d(w748), .e(w427), .x(w426) );
	dmg_aon2222 g804 (.a0(w736), .a1(w486), .b0(w491), .b1(w456), .c0(w102), .c1(w103), .d0(w455), .d1(w105), .x(w944) );
	dmg_aon2222 g805 (.a0(w486), .a1(w485), .b0(w456), .b1(w737), .c0(w103), .c1(w490), .d0(w105), .d1(w106), .x(w772) );
	dmg_aon2222 g806 (.a0(w352), .a1(w838), .b0(w348), .b1(w837), .c0(w357), .c1(w957), .d0(w346), .d1(w345), .x(w773) );
	dmg_aon2222 g807 (.a0(w351), .a1(w352), .b0(w349), .b1(w348), .c0(w358), .c1(w357), .d0(w834), .d1(w346), .x(w946) );
	dmg_aon2222 g808 (.a0(w26), .a1(w391), .b0(w392), .b1(w806), .c0(w98), .c1(w97), .d0(w1), .d1(w864), .x(w786) );
	dmg_aon2222 g809 (.a0(w804), .a1(w26), .b0(w435), .b1(w392), .c0(w99), .c1(w98), .d0(w889), .d1(w1), .x(w2) );
	dmg_aon2222 g810 (.a0(w549), .a1(w550), .b0(w779), .b1(w780), .c0(w481), .c1(w175), .d0(w482), .d1(w655), .x(w654) );
	dmg_or3 g811 (.a(w36), .b(w38), .c(w721), .x(w722) );
	dmg_or3 g812 (.a(w36), .b(w37), .c(w25), .x(w443) );
	dmg_or3 g813 (.a(w36), .b(w445), .c(w23), .x(w22) );
	dmg_or3 g814 (.a(w772), .b(w773), .c(w786), .x(w529) );
	dmg_or3 g815 (.a(w944), .b(w946), .c(w2), .x(w3) );
	dmg_or3 g816 (.a(w36), .b(w783), .c(w784), .x(w436) );
	dmg_or3 g817 (.a(w429), .b(w648), .c(w653), .x(w614) );
	dmg_or3 g818 (.a(w906), .b(w905), .c(w181), .x(w144) );
	dmg_or3 g819 (.a(w36), .b(w40), .c(w193), .x(w194) );
	dmg_or3 g820 (.a(w36), .b(w39), .c(w191), .x(w712) );
	dmg_not3 g821 (.a(w532), .x(w531) );
	dmg_not3 g822 (.a(w423), .x(w422) );
	dmg_not3 g823 (.a(w420), .x(w421) );
	dmg_not3 g824 (.a(w419), .x(w781) );
	dmg_not3 g825 (.a(w6), .x(w5) );
	dmg_not3 g826 (.a(w207), .x(w380) );
	dmg_not3 g827 (.a(w378), .x(w379) );
	dmg_not g828 (.a(w233), .x(w479) );
	dmg_or g829 (.a(w648), .b(w619), .x(w618) );
	dmg_or g830 (.a(w903), .b(w7), .x(w6) );
	dmg_or g831 (.a(w630), .b(w9), .x(w44) );
	dmg_or g832 (.a(w240), .b(w241), .x(w292) );
	dmg_or g833 (.a(w175), .b(w176), .x(w637) );
	dmg_or g834 (.a(w247), .b(w602), .x(w742) );
	dmg_or g835 (.a(w652), .b(w598), .x(w597) );
	dmg_or g836 (.a(w140), .b(w139), .x(w297) );
	dmg_nor g837 (.a(w293), .b(w181), .x(w182) );
	dmg_nand5 g838 (.a(w627), .b(w894), .c(w948), .d(w169), .e(w170), .x(w949) );
	dmg_xor g839 (.a(w245), .b(w246), .x(w616) );
	dmg_xor g840 (.a(w521), .b(w497), .x(w978) );
	dmg_xor g841 (.a(w624), .b(w900), .x(w899) );
	dmg_xor g842 (.a(w815), .b(w814), .x(w901) );
	dmg_xor g843 (.a(w375), .b(w376), .x(w878) );
	dmg_xor g844 (.a(w369), .b(w852), .x(w832) );
	dmg_xor g845 (.a(w286), .b(w856), .x(w417) );
	dmg_xor g846 (.a(w281), .b(w604), .x(w745) );
	dmg_xor g847 (.a(w172), .b(w608), .x(w609) );
	dmg_xor g848 (.a(w361), .b(w879), .x(w746) );
	dmg_xor g849 (.a(w77), .b(w611), .x(w610) );
	dmg_xor g850 (.a(w255), .b(w607), .x(w615) );
	dmg_xor g851 (.a(w252), .b(w750), .x(w418) );
	dmg_xor g852 (.a(w963), .b(w697), .x(w420) );
	dmg_or g853 (.a(w670), .b(w419), .x(w865) );
	dmg_notif1 g854 (.ena(w233), .a(w232), .x(w13) );
	dmg_notif1 g855 (.ena(w210), .a(w562), .x(w48) );
	dmg_notif1 g856 (.ena(w210), .a(w46), .x(w566) );
	dmg_notif1 g857 (.ena(w210), .a(w770), .x(w135) );
	dmg_notif1 g858 (.ena(w210), .a(w858), .x(w126) );
	dmg_notif1 g859 (.ena(w233), .a(w778), .x(w91) );
	dmg_notif1 g860 (.ena(w210), .a(w767), .x(w49) );
	dmg_notif1 g861 (.ena(w210), .a(w766), .x(w60) );
	dmg_notif1 g862 (.ena(w210), .a(w565), .x(w271) );
	dmg_notif1 g863 (.ena(w210), .a(w596), .x(w517) );
	dmg_notif1 g864 (.ena(w210), .a(w209), .x(w65) );
	dmg_notif1 g865 (.ena(w233), .a(w239), .x(w12) );
	dmg_xor g866 (.a(w171), .b(w617), .x(w522) );
	dmg_const g867 (.q0(w14), .q1(w47) );
	dmg_not4 g868 (.a(w904), .x(w630) );
	dmg_not4 g869 (.a(w869), .x(w513) );
	dmg_nor_latch g870 (.s(w754), .r(w637), .q(w636) );
	dmg_nor_latch g871 (.s(w874), .r(w667), .q(w503) );
	dmg_nor_latch g872 (.s(w536), .r(w336), .q(w147) );
	dmg_nor_latch g873 (.s(w150), .r(w151), .q(w75) );
	dmg_nor_latch g874 (.s(w618), .r(w533), .nq(w231) );
	dmg_nor_latch g875 (.s(w523), .r(w618), .q(w524) );
	dmg_nand_latch g876 (.nr(w660), .ns(w143), .q(w764) );
	dmg_nand_latch g877 (.nr(w182), .ns(w823), .q(w183) );
	dmg_or3 g878 (.a(w36), .b(w41), .c(w477), .x(w698) );
	dmg_or3 g879 (.a(w36), .b(w42), .c(w43), .x(w31) );
	dmg_nor g880 (.a(w8), .b(w144), .x(w505) );
	dmg_nor_latch g881 (.s(w8), .r(w7), .q(w9) );
	dmg_dffr_comp g882 (.nr1(w47), .nr2(w47), .d(w311), .ck(w313), .cck(w314), .q(w46) );
	dmg_dffr_comp g883 (.nr1(w47), .nr2(w47), .d(w121), .ck(w313), .cck(w314), .q(w565) );
	dmg_dffr_comp g884 (.nr1(w47), .nr2(w47), .d(w120), .ck(w313), .cck(w314), .q(w562) );
	dmg_dffr_comp g885 (.nr1(w47), .nr2(w47), .d(w554), .ck(w313), .cck(w314), .q(w766) );
	dmg_dffr_comp g886 (.nr1(w47), .nr2(w47), .d(w218), .ck(w313), .cck(w314), .q(w770) );
	dmg_dffr_comp g887 (.nr1(w47), .nr2(w47), .d(w217), .ck(w313), .cck(w314), .q(w858) );
	dmg_dffr_comp g888 (.nr1(w47), .nr2(w47), .d(w553), .ck(w313), .cck(w314), .q(w767) );
	dmg_dffr_comp g889 (.nr1(w47), .nr2(w47), .d(w332), .ck(w313), .cck(w314), .q(w596) );
	dmg_mux g890 (.sel(w122), .d1(w332), .d0(w120), .q(w310) );
	dmg_mux g891 (.sel(w122), .d1(w120), .d0(w332), .q(w886) );
	dmg_mux g892 (.sel(w122), .d1(w554), .d0(w553), .q(w771) );
	dmg_mux g893 (.sel(w122), .d1(w553), .d0(w554), .q(w450) );
	dmg_mux g894 (.sel(w122), .d1(w311), .d0(w121), .q(w459) );
	dmg_mux g895 (.sel(w122), .d1(w121), .d0(w311), .q(w873) );
	dmg_mux g896 (.sel(w122), .d1(w218), .d0(w217), .q(w489) );
	dmg_mux g897 (.sel(w122), .d1(w217), .d0(w218), .q(w448) );
	dmg_nor3 g898 (.a(w533), .b(w898), .c(w144), .x(w143) );
	dmg_nor3 g899 (.a(w667), .b(w469), .c(w470), .x(w463) );
	dmg_nor3 g900 (.a(w534), .b(w535), .c(w851), .x(w823) );
	dmg_nor3 g901 (.a(w620), .b(w500), .c(w659), .x(w915) );
	dmg_nor3 g902 (.a(w178), .b(w179), .c(w176), .x(w177) );
	dmg_nor3 g903 (.a(w598), .b(w526), .c(w227), .x(w226) );
	dmg_nor3 g904 (.a(w868), .b(w598), .c(w205), .x(w204) );
	dmg_nor3 g905 (.a(w441), .b(w440), .c(w439), .x(w438) );
	dmg_nor_latch g906 (.s(w550), .r(w742), .nq(w778) );
	dmg_nand4 g907 (.a(w700), .b(w701), .c(w403), .d(w402), .x(w936) );
	dmg_and4 g908 (.a(w711), .b(w707), .c(w706), .d(w404), .x(w732) );
	dmg_nor3 g909 (.a(w134), .b(w133), .c(w574), .x(w573) );
	dmg_and4 g910 (.a(w77), .b(w281), .c(w255), .d(w252), .x(w544) );
	dmg_nor8 g911 (.a(w77), .b(w281), .c(w255), .d(w252), .e(w286), .f(w245), .g(w361), .h(w172), .x(w425) );
	dmg_and4 g912 (.a(w620), .b(w658), .c(w166), .d(w165), .x(w876) );
	dmg_nand4 g913 (.a(w231), .b(w504), .c(w875), .d(w179), .x(w180) );
	dmg_nor4 g914 (.a(w615), .b(w616), .c(w417), .d(w418), .x(w979) );
	dmg_nor4 g915 (.a(w610), .b(w609), .c(w746), .d(w745), .x(w744) );
	dmg_nand4 g916 (.a(w9), .b(w10), .c(w826), .d(w827), .x(w510) );
endmodule // PPU1

module PPU2 (  cclk, clk6, n_reset2, a, d, n_oamb, oam_bl_pch, oa, n_oam_rd, n_oamb_wr, n_oama_wr, n_oama, CONST0, n_dma_phi, 
	dma_a, dma_run, 
	soc_wr, soc_rd, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, n_ppu_hard_reset, 
	nma, fexx, ff43, ff42, sprite_x_flip, sprite_x_match, bp_sel, ppu_mode3, 
	md, oam_din, v, FF43_D1, FF43_D0, n_ppu_clk, FF43_D2, h, ppu_mode2, vbl, stop_oam_eval, obj_color, vclk2, h_restart, obj_prio_ck, obj_prio, n_ppu_reset, 
	oam_to_vram, n_dma_phi2_latched, FF40_D3, FF40_D2, in_window, 
	FF40_D1, dma_addr_ext, sp_bp_cys, cpu_vram_oam_rd, oam_dma_wr, clk6_delay, oam_mode3_bl_pch, bp_cy, tm_cy, oam_mode3_nrd, ma0, oam_rd_ck, oam_xattr_latch_cck, oam_addr_ck);

	input wire cclk;
	input wire clk6;
	input wire n_reset2;
	input wire [7:0] a;
	inout wire [7:0] d;
	inout wire [7:0] n_oamb;
	output wire oam_bl_pch;
	output wire [7:1] oa; 		// ⚠️ lsb=1
	output wire n_oam_rd;
	output wire n_oamb_wr;
	output wire n_oama_wr;
	inout wire [7:0] n_oama;
	inout wire CONST0;
	input wire n_dma_phi;
	input wire [12:0] dma_a;
	input wire dma_run;
	input wire soc_wr;
	input wire soc_rd;
	output wire ppu_rd;
	output wire ppu_wr;
	output wire ppu_clk;
	input wire vram_to_oam;
	output wire n_ppu_hard_reset;
	inout wire [12:0] nma;
	input wire fexx;
	input wire ff43;
	input wire ff42;
	output wire sprite_x_flip;
	output wire sprite_x_match;
	input wire bp_sel;
	input wire ppu_mode3;
	inout wire [7:0] md;
	output wire FF43_D1;
	output wire FF43_D0;
	output wire n_ppu_clk;
	output wire FF43_D2;
	output wire ppu_mode2;
	input wire vbl;
	output wire stop_oam_eval;
	output wire obj_color;
	input wire vclk2;
	output wire obj_prio;
	input wire n_ppu_reset;
	input wire FF40_D3;
	input wire FF40_D2;
	input wire in_window;
	input wire FF40_D1;
	input wire sp_bp_cys;
	input wire cpu_vram_oam_rd;
	output wire clk6_delay;
	input wire bp_cy;
	input wire tm_cy;
	input wire [7:0] oam_din;
	input wire dma_addr_ext;
	input wire oam_dma_wr;
	input wire obj_prio_ck;
	input wire n_dma_phi2_latched;
	input wire ma0;
	output wire h_restart;
	output wire oam_to_vram;
	input wire oam_mode3_nrd;
	input wire oam_mode3_bl_pch;
	input wire oam_rd_ck;
	input wire oam_xattr_latch_cck;
	input wire oam_addr_ck;

	// H/V
	input wire [7:0] h;
	input wire [7:0] v;

endmodule // PPU2