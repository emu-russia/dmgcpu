
module Decoder2( CLK2, a3, d, w, SeqOut_2 );

	input CLK2;
	input a3;
	input [106:0] d;
	output [40:0] w;
	input SeqOut_2;

endmodule // Decoder2
