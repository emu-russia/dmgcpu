// apu_standalone
// Testing the APU in a spherical vacuum (separate from the other components).
// We just create a APU instance, add all the plugs it needs, and try to get it going.
`timescale 1ns/1ns

module apu_standalone();

endmodule // apu_standalone