module Arbiter (  clk2, n_reset2, cpu_mreq, ext_cs_en, cpu_wr_sync, a, d, cpu_wr, mmio_sel, boot_sel, 
	n_DRV_HIGH_a15, n_INPUT_a15, DRV_LOW_a15, n_cs_topad, CONST0, n_DRV_HIGH_nmwr, n_mwr, DRV_LOW_nmwr, n_DRV_HIGH_nmrd, n_mrd, DRV_LOW_nmrd, n_DRV_HIGH_nmcs, n_mcs, DRV_LOW_nmcs, 
	n_DRV_HIGH_md, n_md_frompad, DRV_LOW_md, n_md_ena_pu, 
	n_DRV_HIGH_d, n_db_frompad, DRV_LOW_d, n_ena_pu_db,
	soc_wr, soc_rd, vram_to_oam, dma_a_15, non_vram_mreq, test_1, n_extdb_to_intdb, n_dblatch_to_intdb, n_intdb_to_extdb, ffxx, n_ppu_hard_reset, ppu_mode3, md, oam_din, n_vram_to_oam, dma_addr_ext, sp_bp_cys, tm_bp_cys, n_sp_bp_mrd, n_tm_bp_cys, arb_fexx_ffxx, cpu_vram_oam_rd);

	input wire clk2;
	input wire n_reset2;
	input wire cpu_mreq;
	input wire ext_cs_en;
	input wire cpu_wr_sync;
	inout wire [15:0] a; 			// ⚠️ a[15] bidir, a[14:0] input
	inout wire [7:0] d;
	input wire cpu_wr;
	output wire mmio_sel;
	output wire boot_sel;
	output wire n_DRV_HIGH_a15;
	input wire n_INPUT_a15;
	output wire DRV_LOW_a15;
	output wire n_cs_topad;
	inout wire CONST0;
	output wire n_DRV_HIGH_nmwr;
	input wire n_mwr;
	output wire DRV_LOW_nmwr;
	output wire n_DRV_HIGH_nmrd;
	input wire n_mrd;
	output wire DRV_LOW_nmrd;
	output wire n_DRV_HIGH_nmcs;
	input wire n_mcs;
	output wire DRV_LOW_nmcs;
	output wire [7:0] n_DRV_HIGH_md;
	input wire [7:0] n_md_frompad;
	output wire [7:0] DRV_LOW_md;
	output wire n_md_ena_pu;
	output wire [7:0] n_DRV_HIGH_d;
	input wire [7:0] n_db_frompad;
	output wire [7:0] DRV_LOW_d;
	input wire n_ena_pu_db;
	input wire soc_wr;
	input wire soc_rd;
	input wire vram_to_oam;
	input wire dma_a_15;
	output wire non_vram_mreq;
	input wire test_1;
	input wire n_extdb_to_intdb;
	input wire n_dblatch_to_intdb;
	input wire n_intdb_to_extdb;
	output wire ffxx;
	input wire n_ppu_hard_reset;
	input wire ppu_mode3;
	inout wire [7:0] md;
	output wire [7:0] oam_din;
	input wire n_vram_to_oam;
	input wire dma_addr_ext;
	input wire sp_bp_cys;
	input wire tm_bp_cys;
	input wire n_tm_bp_cys;
	output wire arb_fexx_ffxx;
	input wire cpu_vram_oam_rd;
	input wire n_sp_bp_mrd;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;

	assign n_DRV_HIGH_d[5] = w1;
	assign w2 = n_INPUT_a15;
	assign DRV_LOW_a15 = w61;
	assign DRV_LOW_d[0] = w62;
	assign n_DRV_HIGH_d[3] = w65;
	assign n_DRV_HIGH_d[0] = w66;
	assign DRV_LOW_d[1] = w228;
	assign n_DRV_HIGH_d[2] = w64;
	assign n_DRV_HIGH_d[1] = w229;
	assign DRV_LOW_d[4] = w63;
	assign w120 = n_db_frompad[5];
	assign n_DRV_HIGH_d[4] = w54;
	assign DRV_LOW_d[3] = w160;
	assign w53 = n_db_frompad[2];
	assign DRV_LOW_d[2] = w161;
	assign n_DRV_HIGH_a15 = w111;
	assign DRV_LOW_d[5] = w110;
	assign w156 = n_db_frompad[1];
	assign w74 = n_db_frompad[3];
	assign w50 = n_db_frompad[0];
	assign w73 = n_db_frompad[4];
	assign DRV_LOW_d[7] = w153;
	assign w152 = n_db_frompad[6];
	assign DRV_LOW_d[6] = w154;
	assign n_DRV_HIGH_d[6] = w221;
	assign w70 = n_db_frompad[7];
	assign n_DRV_HIGH_d[7] = w234;
	assign DRV_LOW_md[0] = w217;
	assign n_DRV_HIGH_md[0] = w218;
	assign DRV_LOW_md[1] = w41;
	assign DRV_LOW_md[6] = w40;
	assign n_md_ena_pu = w42;
	assign n_DRV_HIGH_md[7] = w204;
	assign w211 = n_md_frompad[1];
	assign DRV_LOW_md[7] = w212;
	assign n_DRV_HIGH_md[1] = w203;
	assign w201 = n_md_frompad[7];
	assign w202 = n_md_frompad[2];
	assign n_DRV_HIGH_md[6] = w102;
	assign n_DRV_HIGH_md[2] = w101;
	assign w100 = n_md_frompad[6];
	assign DRV_LOW_md[5] = w37;
	assign n_DRV_HIGH_md[3] = w210;
	assign w209 = n_md_frompad[3];
	assign w208 = n_md_frompad[0];
	assign n_DRV_HIGH_md[5] = w207;
	assign w98 = n_md_frompad[5];
	assign n_DRV_HIGH_md[4] = w105;
	assign DRV_LOW_md[2] = w235;
	assign DRV_LOW_md[4] = w106;
	assign w99 = n_md_frompad[4];
	assign DRV_LOW_md[3] = w213;
	assign w82 = ppu_mode3;
	assign DRV_LOW_nmwr = w83;
	assign n_DRV_HIGH_nmrd = w195;
	assign DRV_LOW_nmrd = w78;
	assign w77 = n_tm_bp_cys;
	assign md[3] = w96;
	assign DRV_LOW_nmcs = w196;
	assign arb_fexx_ffxx = w173;
	assign md[0] = w172;
	assign w149 = tm_bp_cys;
	assign w232 = n_sp_bp_mrd;
	assign n_DRV_HIGH_nmwr = w148;
	assign w144 = n_mwr;
	assign n_DRV_HIGH_nmcs = w145;
	assign md[4] = w56;
	assign md[5] = w35;
	assign md[7] = w34;
	assign w198 = sp_bp_cys;
	assign md[2] = w46;
	assign md[1] = w45;
	assign md[6] = w38;
	assign w88 = n_mrd;
	assign w89 = n_mcs;
	assign w188 = cpu_vram_oam_rd;
	assign w76 = n_vram_to_oam;
	assign oam_din[3] = w75;
	assign oam_din[6] = w151;
	assign w150 = vram_to_oam;
	assign oam_din[0] = w51;
	assign oam_din[2] = w52;
	assign w192 = n_reset2;
	assign oam_din[4] = w72;
	assign oam_din[7] = w71;
	assign w117 = a[6];  		// hand-edited
	assign a[15] = w112;
	assign w9 = n_ppu_hard_reset;
	assign ffxx = w114;
	assign w113 = soc_wr;
	assign oam_din[5] = w119;
	assign w118 = a[4]; 	// hand-edited
	assign w115 = soc_rd;
	assign w131 = a[7]; 	// hand-edited
	assign w132 = a[8]; 	// hand-edited
	assign w133 = a[9]; 	// hand-edited
	assign w134 = a[10]; 	// hand-edited
	assign w135 = a[11]; 	// hand-edited
	assign w136 = a[12]; 	// hand-edited
	assign w126 = a[0]; 	// hand-edited
	assign w127 = a[1]; 	// hand-edited
	assign w128 = a[2]; 	// hand-edited
	assign w129 = a[3]; 	// hand-edited
	assign w130 = a[5]; 	// hand-edited
	assign w138 = a[14]; 	// hand-edited
	assign w137 = a[13]; 	// hand-edited
	assign boot_sel = w225;
	assign w25 = test_1;
	assign w20 = cpu_wr_sync;
	assign w21 = cpu_wr;
	assign d[7] = w5;
	assign non_vram_mreq = w24;
	assign d[0] = w47;
	assign w59 = dma_a_15;
	assign d[6] = w31;
	assign d[5] = w28;
	assign w29 = dma_addr_ext;
	assign w68 = n_extdb_to_intdb;
	assign w159 = n_dblatch_to_intdb;
	assign d[4] = w55;
	assign w30 = n_intdb_to_extdb;
	assign CONST0 = w165;
	assign d[3] = w27;
	assign mmio_sel = w178;
	assign w177 = cpu_mreq;
	assign d[2] = w108;
	assign d[1] = w122;
	assign n_cs_topad = w184;
	assign w93 = clk2;
	assign w92 = ext_cs_en;
	assign oam_din[1] = w233;
	assign w48 = n_ena_pu_db;

	// Instances

	dmg_nand g1 (.a(w28), .b(w48), .x(w1) );
	dmg_nand g2 (.a(w27), .b(w48), .x(w65) );
	dmg_nand g3 (.a(w108), .b(w48), .x(w64) );
	dmg_nand g4 (.a(w47), .b(w48), .x(w66) );
	dmg_nand g5 (.a(w122), .b(w48), .x(w229) );
	dmg_nand g6 (.a(w5), .b(w48), .x(w234) );
	dmg_nand g7 (.a(w31), .b(w48), .x(w221) );
	dmg_nand g8 (.a(w15), .b(w16), .x(w81) );
	dmg_nand g9 (.a(w226), .b(w141), .x(w143) );
	dmg_nand g10 (.a(w92), .b(w57), .x(w58) );
	dmg_not g11 (.a(w53), .x(w67) );
	dmg_not g12 (.a(w156), .x(w157) );
	dmg_not g13 (.a(w2), .x(w3) );
	dmg_not g14 (.a(w120), .x(w121) );
	dmg_not g15 (.a(w25), .x(w4) );
	dmg_not g16 (.a(w70), .x(w69) );
	dmg_not g17 (.a(w32), .x(w33) );
	dmg_not g18 (.a(w46), .x(w107) );
	dmg_not g19 (.a(w45), .x(w123) );
	dmg_not g20 (.a(w96), .x(w95) );
	dmg_not g21 (.a(w38), .x(w183) );
	dmg_not g22 (.a(w35), .x(w182) );
	dmg_not g23 (.a(w172), .x(w230) );
	dmg_not g24 (.a(w12), .x(w43) );
	dmg_not g25 (.a(w14), .x(w13) );
	dmg_not g26 (.a(w11), .x(w14) );
	dmg_not g27 (.a(w15), .x(w140) );
	dmg_not g28 (.a(w50), .x(w51) );
	dmg_not g29 (.a(w139), .x(w173) );
	dmg_not g30 (.a(w82), .x(w16) );
	dmg_not g31 (.a(w86), .x(w85) );
	dmg_and g32 (.a(w177), .b(w176), .x(w24) );
	dmg_and g33 (.a(w38), .b(w33), .x(w103) );
	dmg_and g34 (.a(w45), .b(w33), .x(w44) );
	dmg_and g35 (.a(w35), .b(w33), .x(w220) );
	dmg_and g36 (.a(w46), .b(w33), .x(w215) );
	dmg_and g37 (.a(w172), .b(w33), .x(w219) );
	dmg_and g38 (.a(w96), .b(w33), .x(w97) );
	dmg_and g39 (.a(w56), .b(w33), .x(w206) );
	dmg_and g40 (.a(w34), .b(w33), .x(w205) );
	dmg_and g41 (.a(w112), .b(w23), .x(w22) );
	dmg_and g42 (.a(w141), .b(w140), .x(w11) );
	dmg_and g43 (.a(w17), .b(w16), .x(w141) );
	dmg_and g44 (.a(w80), .b(w85), .x(w194) );
	dmg_and g45 (.a(w11), .b(w13), .x(w231) );
	dmg_nor g46 (.a(w30), .b(w47), .x(w62) );
	dmg_nor g47 (.a(w30), .b(w55), .x(w63) );
	dmg_nor g48 (.a(w30), .b(w122), .x(w228) );
	dmg_nor g49 (.a(w60), .b(w25), .x(w61) );
	dmg_nor g50 (.a(w30), .b(w5), .x(w153) );
	dmg_nor g51 (.a(w30), .b(w31), .x(w154) );
	dmg_nor g52 (.a(w189), .b(w139), .x(w114) );
	dmg_nor g53 (.a(w112), .b(w225), .x(w57) );
	dmg_nor g54 (.a(w30), .b(w108), .x(w161) );
	dmg_nor g55 (.a(w30), .b(w27), .x(w160) );
	dmg_nor g56 (.a(w30), .b(w28), .x(w110) );
	dmg_nor g57 (.a(w25), .b(w93), .x(w94) );
	dmg_nor g58 (.a(w178), .b(w24), .x(w23) );
	dmg_nand g59 (.a(w141), .b(w188), .x(w193) );
	dmg_not2 g60 (.a(w197), .x(w196) );
	dmg_not2 g61 (.a(w194), .x(w195) );
	dmg_not2 g62 (.a(w84), .x(w83) );
	dmg_not2 g63 (.a(w79), .x(w78) );
	dmg_not2 g64 (.a(w214), .x(w235) );
	dmg_not2 g65 (.a(w181), .x(w106) );
	dmg_not2 g66 (.a(w199), .x(w212) );
	dmg_not2 g67 (.a(w200), .x(w213) );
	dmg_not2 g68 (.a(w205), .x(w204) );
	dmg_not2 g69 (.a(w97), .x(w210) );
	dmg_not2 g70 (.a(w215), .x(w101) );
	dmg_not2 g71 (.a(w44), .x(w203) );
	dmg_not2 g72 (.a(w36), .x(w37) );
	dmg_not2 g73 (.a(w43), .x(w42) );
	dmg_not2 g74 (.a(w104), .x(w41) );
	dmg_not2 g75 (.a(w103), .x(w102) );
	dmg_not2 g76 (.a(w206), .x(w105) );
	dmg_not2 g77 (.a(w39), .x(w40) );
	dmg_not2 g78 (.a(w220), .x(w207) );
	dmg_not2 g79 (.a(w219), .x(w218) );
	dmg_not2 g80 (.a(w216), .x(w217) );
	dmg_not2 g81 (.a(w94), .x(w49) );
	dmg_not2 g82 (.a(w147), .x(w148) );
	dmg_not2 g83 (.a(w146), .x(w145) );
	dmg_not g84 (.a(w132), .x(w189) );
	dmg_nand g85 (.a(w55), .b(w48), .x(w54) );
	dmg_notif0 g86 (.n_ena(w159), .a(w155), .x(w122) );
	dmg_notif0 g87 (.n_ena(w159), .a(w162), .x(w47) );
	dmg_notif0 g88 (.n_ena(w159), .a(w163), .x(w108) );
	dmg_notif1 g89 (.ena(w43), .a(w211), .x(w45) );
	dmg_notif1 g90 (.ena(w43), .a(w100), .x(w38) );
	dmg_notif1 g91 (.ena(w43), .a(w202), .x(w46) );
	dmg_notif1 g92 (.ena(w43), .a(w98), .x(w35) );
	dmg_notif1 g93 (.ena(w43), .a(w209), .x(w96) );
	dmg_notif1 g94 (.ena(w43), .a(w208), .x(w172) );
	dmg_notif1 g95 (.ena(w43), .a(w201), .x(w34) );
	dmg_notif1 g96 (.ena(w43), .a(w99), .x(w56) );
	dmg_notif1 g97 (.ena(w7), .a(w107), .x(w108) );
	dmg_notif1 g98 (.ena(w7), .a(w123), .x(w122) );
	dmg_notif1 g99 (.ena(w7), .a(w95), .x(w27) );
	dmg_notif1 g100 (.ena(w7), .a(w183), .x(w31) );
	dmg_notif1 g101 (.ena(w7), .a(w182), .x(w28) );
	dmg_notif1 g102 (.ena(w7), .a(w230), .x(w47) );
	dmg_notif1 g103 (.ena(w190), .a(w171), .x(w47) );
	dmg_notif0 g104 (.n_ena(w159), .a(w222), .x(w28) );
	dmg_notif0 g105 (.n_ena(w159), .a(w164), .x(w31) );
	dmg_notif0 g106 (.n_ena(w159), .a(w158), .x(w27) );
	dmg_notif0 g107 (.n_ena(w159), .a(w223), .x(w55) );
	dmg_notif0 g108 (.n_ena(w159), .a(w166), .x(w5) );
	dmg_notif1 g109 (.ena(w7), .a(w124), .x(w55) );
	dmg_bufif0 g110 (.a0(w28), .n_ena(w32), .a1(w28), .x(w35) );
	dmg_bufif0 g111 (.a0(w69), .n_ena(w68), .a1(w69), .x(w5) );
	dmg_bufif0 g112 (.a0(w67), .n_ena(w68), .a1(w67), .x(w108) );
	dmg_bufif0 g113 (.a0(w157), .n_ena(w68), .a1(w157), .x(w122) );
	dmg_bufif0 g114 (.a0(w121), .n_ena(w68), .a1(w121), .x(w28) );
	dmg_bufif0 g115 (.a0(w26), .n_ena(w49), .a1(w26), .x(w122) );
	dmg_bufif0 g116 (.a0(w26), .n_ena(w49), .a1(w26), .x(w108) );
	dmg_bufif0 g117 (.a0(w3), .n_ena(w4), .a1(w3), .x(w112) );
	dmg_bufif0 g118 (.a0(w5), .n_ena(w32), .a1(w5), .x(w34) );
	dmg_bufif0 g119 (.a0(w27), .n_ena(w32), .a1(w27), .x(w96) );
	dmg_bufif0 g120 (.a0(w55), .n_ena(w32), .a1(w55), .x(w56) );
	dmg_bufif0 g121 (.a0(w47), .n_ena(w32), .a1(w47), .x(w172) );
	dmg_bufif0 g122 (.a0(w108), .n_ena(w32), .a1(w108), .x(w46) );
	dmg_bufif0 g123 (.a0(w31), .n_ena(w32), .a1(w31), .x(w38) );
	dmg_bufif0 g124 (.a0(w122), .n_ena(w32), .a1(w122), .x(w45) );
	dmg_bufif0 g125 (.a0(w186), .n_ena(w68), .a1(w186), .x(w47) );
	dmg_bufif0 g126 (.a0(w185), .n_ena(w68), .a1(w185), .x(w31) );
	dmg_bufif0 g127 (.a0(w26), .n_ena(w49), .a1(w26), .x(w5) );
	dmg_bufif0 g128 (.a0(w26), .n_ena(w49), .a1(w26), .x(w31) );
	dmg_bufif0 g129 (.a0(w26), .n_ena(w49), .a1(w26), .x(w47) );
	dmg_bufif0 g130 (.a0(w26), .n_ena(w49), .a1(w26), .x(w27) );
	dmg_bufif0 g131 (.a0(w26), .n_ena(w49), .a1(w26), .x(w28) );
	dmg_bufif0 g132 (.a0(w26), .n_ena(w49), .a1(w26), .x(w55) );
	dmg_bufif0 g133 (.a0(w227), .n_ena(w68), .a1(w227), .x(w55) );
	dmg_bufif0 g134 (.a0(w109), .n_ena(w68), .a1(w109), .x(w27) );
	dmg_latch g135 (.ena(w159), .d(w156), .q(w155) );
	dmg_latch g136 (.ena(w159), .d(w53), .q(w163) );
	dmg_latch g137 (.ena(w159), .d(w152), .q(w164) );
	dmg_latch g138 (.ena(w159), .d(w70), .q(w166) );
	dmg_latch g139 (.ena(w159), .d(w120), .q(w222) );
	dmg_latch g140 (.ena(w159), .d(w73), .q(w223) );
	dmg_latch g141 (.ena(w159), .d(w50), .q(w162) );
	dmg_latch g142 (.ena(w159), .d(w74), .q(w158) );
	dmg_notif1 g143 (.ena(w7), .a(w6), .x(w5) );
	dmg_or g144 (.a(w86), .b(w80), .x(w79) );
	dmg_or g145 (.a(w13), .b(w11), .x(w12) );
	dmg_or g146 (.a(w32), .b(w46), .x(w214) );
	dmg_or g147 (.a(w32), .b(w45), .x(w104) );
	dmg_or g148 (.a(w32), .b(w38), .x(w39) );
	dmg_or g149 (.a(w32), .b(w35), .x(w36) );
	dmg_or g150 (.a(w32), .b(w172), .x(w216) );
	dmg_or g151 (.a(w32), .b(w96), .x(w200) );
	dmg_or g152 (.a(w32), .b(w34), .x(w199) );
	dmg_or g153 (.a(w32), .b(w56), .x(w181) );
	dmg_or g154 (.a(w47), .b(w170), .x(w191) );
	dmg_or g155 (.a(w86), .b(w143), .x(w84) );
	dmg_or g156 (.a(w86), .b(w142), .x(w197) );
	dmg_nand g157 (.a(w60), .b(w4), .x(w111) );
	dmg_nand g158 (.a(w22), .b(w21), .x(w174) );
	dmg_mux g159 (.sel(w29), .d1(w59), .d0(w58), .q(w60) );
	dmg_mux g160 (.sel(w29), .d1(w59), .d0(w167), .q(w184) );
	dmg_mux g161 (.sel(w86), .d1(w90), .d0(w91), .q(w17) );
	dmg_mux g162 (.sel(w86), .d1(w18), .d0(w19), .q(w226) );
	dmg_mux g163 (.sel(w86), .d1(w87), .d0(w174), .q(w15) );
	dmg_not3 g164 (.a(w231), .x(w32) );
	dmg_and4 g165 (.a(w81), .b(w232), .c(w77), .d(w76), .x(w80) );
	dmg_dffr g166 (.clk(w8), .nr1(w9), .nr2(w9), .d(w10), .nq(w10) );
	dmg_dffr g167 (.clk(w187), .nr1(w192), .nr2(w192), .d(w191), .nq(w171), .q(w170) );
	dmg_or3 g168 (.a(w137), .b(w138), .c(w224), .x(w176) );
	dmg_and3 g169 (.a(w175), .b(w92), .c(w139), .x(w167) );
	dmg_and3 g170 (.a(w137), .b(w180), .c(w112), .x(w179) );
	dmg_nand4 g171 (.a(w125), .b(w116), .c(w114), .d(w113), .x(w187) );
	dmg_and4 g172 (.a(w115), .b(w114), .c(w116), .d(w125), .x(w190) );
	dmg_nor8 g173 (.a(w112), .b(w138), .c(w137), .d(w136), .e(w135), .f(w134), .g(w133), .h(w132), .x(w168) );
	dmg_nand7 g174 (.a(w112), .b(w138), .c(w137), .d(w136), .e(w135), .f(w133), .g(w133), .x(w139) );
	dmg_nor6 g175 (.a(w131), .b(w130), .c(w129), .d(w128), .e(w127), .f(w126), .x(w125) );
	dmg_nor4 g176 (.a(w149), .b(w150), .c(w198), .d(w141), .x(w142) );
	dmg_const g177 (.q0(w165), .q1(w26) );
	dmg_aon g178 (.a0(w112), .a1(w138), .b(w179), .x(w175) );
	dmg_not g179 (.a(w144), .x(w18) );
	dmg_not g180 (.a(w53), .x(w52) );
	dmg_not g181 (.a(w25), .x(w8) );
	dmg_not g182 (.a(w193), .x(w7) );
	dmg_not g183 (.a(w73), .x(w72) );
	dmg_not g184 (.a(w56), .x(w124) );
	dmg_not g185 (.a(w120), .x(w119) );
	dmg_not g186 (.a(w70), .x(w71) );
	dmg_not g187 (.a(w34), .x(w6) );
	dmg_not g188 (.a(w138), .x(w180) );
	dmg_not g189 (.a(w139), .x(w178) );
	dmg_not g190 (.a(w112), .x(w224) );
	dmg_not g191 (.a(w152), .x(w185) );
	dmg_not g192 (.a(w74), .x(w109) );
	dmg_not g193 (.a(w73), .x(w227) );
	dmg_not g194 (.a(w156), .x(w233) );
	dmg_not g195 (.a(w170), .x(w169) );
	dmg_not g196 (.a(w50), .x(w186) );
	dmg_not g197 (.a(w88), .x(w87) );
	dmg_not g198 (.a(w152), .x(w151) );
	dmg_not g199 (.a(w89), .x(w90) );
	dmg_not g200 (.a(w74), .x(w75) );
	dmg_and g201 (.a(w142), .b(w85), .x(w146) );
	dmg_and g202 (.a(w143), .b(w85), .x(w147) );
	dmg_and g203 (.a(w25), .b(w10), .x(w86) );
	dmg_and g204 (.a(w118), .b(w117), .x(w116) );
	dmg_and g205 (.a(w169), .b(w168), .x(w225) );
	dmg_and g206 (.a(w22), .b(w20), .x(w19) );
	dmg_and g207 (.a(w22), .b(w92), .x(w91) );
endmodule // Arbiter