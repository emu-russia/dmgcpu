module PPU1 (  a, d, n_ma, n_lcd_ld1, n_lcd_ld0, n_lcd_cpg, n_lcd_cp, n_lcd_st, n_lcd_cpl, n_lcd_fr, n_lcd_s, CONST0, n_dma_phi, ppu_rd, ppu_wr, ppu_clk, vram_to_oam, ffxx, n_ppu_hard_reset, ff46, 
	nma, fexx, ff43, ff42, sprite_x_flip, sprite_x_match, bp_sel, ppu_mode3, 
	md, v, FF43_D1, FF43_D0, n_ppu_clk, FF43_D2, h, ppu_mode2, vbl, stop_oam_eval, obj_color, vclk2, h_restart, obj_prio_ck, obj_prio, n_ppu_reset, n_dma_phi2_latched, FF40_D3, FF40_D2, in_window, 
	FF40_D1, sp_bp_cys, tm_bp_cys, n_sp_bp_mrd, n_tm_bp_cys, arb_fexx_ffxx, ppu_int_stat, ppu_int_vbl, oam_mode3_bl_pch, bp_cy, tm_cy, oam_mode3_nrd, ppu1_ma0, oam_rd_ck, oam_xattr_latch_cck, oam_addr_ck);

	input wire [12:0] a;
	inout wire [7:0] d;
	output wire [12:0] n_ma;
	output wire n_lcd_ld1;
	output wire n_lcd_ld0;
	output wire n_lcd_cpg;
	output wire n_lcd_cp;
	output wire n_lcd_st;
	output wire n_lcd_cpl;
	output wire n_lcd_fr;
	output wire n_lcd_s;
	inout wire CONST0;
	input wire n_dma_phi;
	input wire ppu_rd;
	input wire ppu_wr;
	input wire ppu_clk;
	input wire vram_to_oam;
	input wire ffxx;
	input wire n_ppu_hard_reset;
	output wire ff46;
	inout wire [12:0] nma;
	output wire fexx;
	output wire ff43;
	output wire ff42;
	input wire sprite_x_flip;
	input wire sprite_x_match;
	output wire bp_sel;
	output wire ppu_mode3;
	inout wire [7:0] md;
	input wire FF43_D1;
	input wire FF43_D0;
	input wire n_ppu_clk;
	input wire FF43_D2;
	input wire ppu_mode2;
	output wire vbl;
	input wire stop_oam_eval;
	input wire obj_color;
	output wire vclk2;
	input wire obj_prio;
	output wire n_ppu_reset;
	output wire FF40_D3;
	output wire FF40_D2;
	output wire in_window;
	output wire FF40_D1;
	output wire sp_bp_cys;
	output wire tm_bp_cys;
	output wire n_tm_bp_cys;
	input wire arb_fexx_ffxx;
	output wire ppu_int_stat;
	output wire ppu_int_vbl;
	output wire bp_cy;
	output wire tm_cy;
	input wire h_restart;
	output wire obj_prio_ck;
	output wire n_dma_phi2_latched;
	output wire ppu1_ma0;
	output wire n_sp_bp_mrd; 		// to arb

	output wire oam_mode3_nrd;  		// is low when OAM is read during MODE3 (pixel transfer stage)
	output wire oam_mode3_bl_pch;
	// @msinger: I guess you already noticed yourself that XUJY(oam_mode3_bl_pch) is the same as XUJA(oam_mode3_nrd), but it is low for a little bit longer.
	// I don't know why it is longer, but it seems to be used to control the OAM bitline precharging during MODE3. It disables the precharging temporarily so that the read access can be performed.   (#328)

	// OAM Clocks
	output wire oam_rd_ck;
	output wire oam_xattr_latch_cck;
	output wire oam_addr_ck;

	// H/V

	output wire [7:0] h;
	output wire [7:0] v;

	// Wires

	wire w1;
	wire w2;
	wire w3;
	wire w4;
	wire w5;
	wire w6;
	wire w7;
	wire w8;
	wire w9;
	wire w10;
	wire w11;
	wire w12;
	wire w13;
	wire w14;
	wire w15;
	wire w16;
	wire w17;
	wire w18;
	wire w19;
	wire w20;
	wire w21;
	wire w22;
	wire w23;
	wire w24;
	wire w25;
	wire w26;
	wire w27;
	wire w28;
	wire w29;
	wire w30;
	wire w31;
	wire w32;
	wire w33;
	wire w34;
	wire w35;
	wire w36;
	wire w37;
	wire w38;
	wire w39;
	wire w40;
	wire w41;
	wire w42;
	wire w43;
	wire w44;
	wire w45;
	wire w46;
	wire w47;
	wire w48;
	wire w49;
	wire w50;
	wire w51;
	wire w52;
	wire w53;
	wire w54;
	wire w55;
	wire w56;
	wire w57;
	wire w58;
	wire w59;
	wire w60;
	wire w61;
	wire w62;
	wire w63;
	wire w64;
	wire w65;
	wire w66;
	wire w67;
	wire w68;
	wire w69;
	wire w70;
	wire w71;
	wire w72;
	wire w73;
	wire w74;
	wire w75;
	wire w76;
	wire w77;
	wire w78;
	wire w79;
	wire w80;
	wire w81;
	wire w82;
	wire w83;
	wire w84;
	wire w85;
	wire w86;
	wire w87;
	wire w88;
	wire w89;
	wire w90;
	wire w91;
	wire w92;
	wire w93;
	wire w94;
	wire w95;
	wire w96;
	wire w97;
	wire w98;
	wire w99;
	wire w100;
	wire w101;
	wire w102;
	wire w103;
	wire w104;
	wire w105;
	wire w106;
	wire w107;
	wire w108;
	wire w109;
	wire w110;
	wire w111;
	wire w112;
	wire w113;
	wire w114;
	wire w115;
	wire w116;
	wire w117;
	wire w118;
	wire w119;
	wire w120;
	wire w121;
	wire w122;
	wire w123;
	wire w124;
	wire w125;
	wire w126;
	wire w127;
	wire w128;
	wire w129;
	wire w130;
	wire w131;
	wire w132;
	wire w133;
	wire w134;
	wire w135;
	wire w136;
	wire w137;
	wire w138;
	wire w139;
	wire w140;
	wire w141;
	wire w142;
	wire w143;
	wire w144;
	wire w145;
	wire w146;
	wire w147;
	wire w148;
	wire w149;
	wire w150;
	wire w151;
	wire w152;
	wire w153;
	wire w154;
	wire w155;
	wire w156;
	wire w157;
	wire w158;
	wire w159;
	wire w160;
	wire w161;
	wire w162;
	wire w163;
	wire w164;
	wire w165;
	wire w166;
	wire w167;
	wire w168;
	wire w169;
	wire w170;
	wire w171;
	wire w172;
	wire w173;
	wire w174;
	wire w175;
	wire w176;
	wire w177;
	wire w178;
	wire w179;
	wire w180;
	wire w181;
	wire w182;
	wire w183;
	wire w184;
	wire w185;
	wire w186;
	wire w187;
	wire w188;
	wire w189;
	wire w190;
	wire w191;
	wire w192;
	wire w193;
	wire w194;
	wire w195;
	wire w196;
	wire w197;
	wire w198;
	wire w199;
	wire w200;
	wire w201;
	wire w202;
	wire w203;
	wire w204;
	wire w205;
	wire w206;
	wire w207;
	wire w208;
	wire w209;
	wire w210;
	wire w211;
	wire w212;
	wire w213;
	wire w214;
	wire w215;
	wire w216;
	wire w217;
	wire w218;
	wire w219;
	wire w220;
	wire w221;
	wire w222;
	wire w223;
	wire w224;
	wire w225;
	wire w226;
	wire w227;
	wire w228;
	wire w229;
	wire w230;
	wire w231;
	wire w232;
	wire w233;
	wire w234;
	wire w235;
	wire w236;
	wire w237;
	wire w238;
	wire w239;
	wire w240;
	wire w241;
	wire w242;
	wire w243;
	wire w244;
	wire w245;
	wire w246;
	wire w247;
	wire w248;
	wire w249;
	wire w250;
	wire w251;
	wire w252;
	wire w253;
	wire w254;
	wire w255;
	wire w256;
	wire w257;
	wire w258;
	wire w259;
	wire w260;
	wire w261;
	wire w262;
	wire w263;
	wire w264;
	wire w265;
	wire w266;
	wire w267;
	wire w268;
	wire w269;
	wire w270;
	wire w271;
	wire w272;
	wire w273;
	wire w274;
	wire w275;
	wire w276;
	wire w277;
	wire w278;
	wire w279;
	wire w280;
	wire w281;
	wire w282;
	wire w283;
	wire w284;
	wire w285;
	wire w286;
	wire w287;
	wire w288;
	wire w289;
	wire w290;
	wire w291;
	wire w292;
	wire w293;
	wire w294;
	wire w295;
	wire w296;
	wire w297;
	wire w298;
	wire w299;
	wire w300;
	wire w301;
	wire w302;
	wire w303;
	wire w304;
	wire w305;
	wire w306;
	wire w307;
	wire w308;
	wire w309;
	wire w310;
	wire w311;
	wire w312;
	wire w313;
	wire w314;
	wire w315;
	wire w316;
	wire w317;
	wire w318;
	wire w319;
	wire w320;
	wire w321;
	wire w322;
	wire w323;
	wire w324;
	wire w325;
	wire w326;
	wire w327;
	wire w328;
	wire w329;
	wire w330;
	wire w331;
	wire w332;
	wire w333;
	wire w334;
	wire w335;
	wire w336;
	wire w337;
	wire w338;
	wire w339;
	wire w340;
	wire w341;
	wire w342;
	wire w343;
	wire w344;
	wire w345;
	wire w346;
	wire w347;
	wire w348;
	wire w349;
	wire w350;
	wire w351;
	wire w352;
	wire w353;
	wire w354;
	wire w355;
	wire w356;
	wire w357;
	wire w358;
	wire w359;
	wire w360;
	wire w361;
	wire w362;
	wire w363;
	wire w364;
	wire w365;
	wire w366;
	wire w367;
	wire w368;
	wire w369;
	wire w370;
	wire w371;
	wire w372;
	wire w373;
	wire w374;
	wire w375;
	wire w376;
	wire w377;
	wire w378;
	wire w379;
	wire w380;
	wire w381;
	wire w382;
	wire w383;
	wire w384;
	wire w385;
	wire w386;
	wire w387;
	wire w388;
	wire w389;
	wire w390;
	wire w391;
	wire w392;
	wire w393;
	wire w394;
	wire w395;
	wire w396;
	wire w397;
	wire w398;
	wire w399;
	wire w400;
	wire w401;
	wire w402;
	wire w403;
	wire w404;
	wire w405;
	wire w406;
	wire w407;
	wire w408;
	wire w409;
	wire w410;
	wire w411;
	wire w412;
	wire w413;
	wire w414;
	wire w415;
	wire w416;
	wire w417;
	wire w418;
	wire w419;
	wire w420;
	wire w421;
	wire w422;
	wire w423;
	wire w424;
	wire w425;
	wire w426;
	wire w427;
	wire w428;
	wire w429;
	wire w430;
	wire w431;
	wire w432;
	wire w433;
	wire w434;
	wire w435;
	wire w436;
	wire w437;
	wire w438;
	wire w439;
	wire w440;
	wire w441;
	wire w442;
	wire w443;
	wire w444;
	wire w445;
	wire w446;
	wire w447;
	wire w448;
	wire w449;
	wire w450;
	wire w451;
	wire w452;
	wire w453;
	wire w454;
	wire w455;
	wire w456;
	wire w457;
	wire w458;
	wire w459;
	wire w460;
	wire w461;
	wire w462;
	wire w463;
	wire w464;
	wire w465;
	wire w466;
	wire w467;
	wire w468;
	wire w469;
	wire w470;
	wire w471;
	wire w472;
	wire w473;
	wire w474;
	wire w475;
	wire w476;
	wire w477;
	wire w478;
	wire w479;
	wire w480;
	wire w481;
	wire w482;
	wire w483;
	wire w484;
	wire w485;
	wire w486;
	wire w487;
	wire w488;
	wire w489;
	wire w490;
	wire w491;
	wire w492;
	wire w493;
	wire w494;
	wire w495;
	wire w496;
	wire w497;
	wire w498;
	wire w499;
	wire w500;
	wire w501;
	wire w502;
	wire w503;
	wire w504;
	wire w505;
	wire w506;
	wire w507;
	wire w508;
	wire w509;
	wire w510;
	wire w511;
	wire w512;
	wire w513;
	wire w514;
	wire w515;
	wire w516;
	wire w517;
	wire w518;
	wire w519;
	wire w520;
	wire w521;
	wire w522;
	wire w523;
	wire w524;
	wire w525;
	wire w526;
	wire w527;
	wire w528;
	wire w529;
	wire w530;
	wire w531;
	wire w532;
	wire w533;
	wire w534;
	wire w535;
	wire w536;
	wire w537;
	wire w538;
	wire w539;
	wire w540;
	wire w541;
	wire w542;
	wire w543;
	wire w544;
	wire w545;
	wire w546;
	wire w547;
	wire w548;
	wire w549;
	wire w550;
	wire w551;
	wire w552;
	wire w553;
	wire w554;
	wire w555;
	wire w556;
	wire w557;
	wire w558;
	wire w559;
	wire w560;
	wire w561;
	wire w562;
	wire w563;
	wire w564;
	wire w565;
	wire w566;
	wire w567;
	wire w568;
	wire w569;
	wire w570;
	wire w571;
	wire w572;
	wire w573;
	wire w574;
	wire w575;
	wire w576;
	wire w577;
	wire w578;
	wire w579;
	wire w580;
	wire w581;
	wire w582;
	wire w583;
	wire w584;
	wire w585;
	wire w586;
	wire w587;
	wire w588;
	wire w589;
	wire w590;
	wire w591;
	wire w592;
	wire w593;
	wire w594;
	wire w595;
	wire w596;
	wire w597;
	wire w598;
	wire w599;
	wire w600;
	wire w601;
	wire w602;
	wire w603;
	wire w604;
	wire w605;
	wire w606;
	wire w607;
	wire w608;
	wire w609;
	wire w610;
	wire w611;
	wire w612;
	wire w613;
	wire w614;
	wire w615;
	wire w616;
	wire w617;
	wire w618;
	wire w619;
	wire w620;
	wire w621;
	wire w622;
	wire w623;
	wire w624;
	wire w625;
	wire w626;
	wire w627;
	wire w628;
	wire w629;
	wire w630;
	wire w631;
	wire w632;
	wire w633;
	wire w634;
	wire w635;
	wire w636;
	wire w637;
	wire w638;
	wire w639;
	wire w640;
	wire w641;
	wire w642;
	wire w643;
	wire w644;
	wire w645;
	wire w646;
	wire w647;
	wire w648;
	wire w649;
	wire w650;
	wire w651;
	wire w652;
	wire w653;
	wire w654;
	wire w655;
	wire w656;
	wire w657;
	wire w658;
	wire w659;
	wire w660;
	wire w661;
	wire w662;
	wire w663;
	wire w664;
	wire w665;
	wire w666;
	wire w667;
	wire w668;
	wire w669;
	wire w670;
	wire w671;
	wire w672;
	wire w673;
	wire w674;
	wire w675;
	wire w676;
	wire w677;
	wire w678;
	wire w679;
	wire w680;
	wire w681;
	wire w682;
	wire w683;
	wire w684;
	wire w685;
	wire w686;
	wire w687;
	wire w688;
	wire w689;
	wire w690;
	wire w691;
	wire w692;
	wire w693;
	wire w694;
	wire w695;
	wire w696;
	wire w697;
	wire w698;
	wire w699;
	wire w700;
	wire w701;
	wire w702;
	wire w703;
	wire w704;
	wire w705;
	wire w706;
	wire w707;
	wire w708;
	wire w709;
	wire w710;
	wire w711;
	wire w712;
	wire w713;
	wire w714;
	wire w715;
	wire w716;
	wire w717;
	wire w718;
	wire w719;
	wire w720;
	wire w721;
	wire w722;
	wire w723;
	wire w724;
	wire w725;
	wire w726;
	wire w727;
	wire w728;
	wire w729;
	wire w730;
	wire w731;
	wire w732;
	wire w733;
	wire w734;
	wire w735;
	wire w736;
	wire w737;
	wire w738;
	wire w739;
	wire w740;
	wire w741;
	wire w742;
	wire w743;
	wire w744;
	wire w745;
	wire w746;
	wire w747;
	wire w748;
	wire w749;
	wire w750;
	wire w751;
	wire w752;
	wire w753;
	wire w754;
	wire w755;
	wire w756;
	wire w757;
	wire w758;
	wire w759;
	wire w760;
	wire w761;
	wire w762;
	wire w763;
	wire w764;
	wire w765;
	wire w766;
	wire w767;
	wire w768;
	wire w769;
	wire w770;
	wire w771;
	wire w772;
	wire w773;
	wire w774;
	wire w775;
	wire w776;
	wire w777;
	wire w778;
	wire w779;
	wire w780;
	wire w781;
	wire w782;
	wire w783;
	wire w784;
	wire w785;
	wire w786;
	wire w787;
	wire w788;
	wire w789;
	wire w790;
	wire w791;
	wire w792;
	wire w793;
	wire w794;
	wire w795;
	wire w796;
	wire w797;
	wire w798;
	wire w799;
	wire w800;
	wire w801;
	wire w802;
	wire w803;
	wire w804;
	wire w805;
	wire w806;
	wire w807;
	wire w808;
	wire w809;
	wire w810;
	wire w811;
	wire w812;
	wire w813;
	wire w814;
	wire w815;
	wire w816;
	wire w817;
	wire w818;
	wire w819;
	wire w820;
	wire w821;
	wire w822;
	wire w823;
	wire w824;
	wire w825;
	wire w826;
	wire w827;
	wire w828;
	wire w829;
	wire w830;
	wire w831;
	wire w832;
	wire w833;
	wire w834;
	wire w835;
	wire w836;
	wire w837;
	wire w838;
	wire w839;
	wire w840;
	wire w841;
	wire w842;
	wire w843;
	wire w844;
	wire w845;
	wire w846;
	wire w847;
	wire w848;
	wire w849;
	wire w850;
	wire w851;
	wire w852;
	wire w853;
	wire w854;
	wire w855;
	wire w856;
	wire w857;
	wire w858;
	wire w859;
	wire w860;
	wire w861;
	wire w862;
	wire w863;
	wire w864;
	wire w865;
	wire w866;
	wire w867;
	wire w868;
	wire w869;
	wire w870;
	wire w871;
	wire w872;
	wire w873;
	wire w874;
	wire w875;
	wire w876;
	wire w877;
	wire w878;
	wire w879;
	wire w880;
	wire w881;
	wire w882;
	wire w883;
	wire w884;
	wire w885;
	wire w886;
	wire w887;
	wire w888;
	wire w889;
	wire w890;
	wire w891;
	wire w892;
	wire w893;
	wire w894;
	wire w895;
	wire w896;
	wire w897;
	wire w898;
	wire w899;
	wire w900;
	wire w901;
	wire w902;
	wire w903;
	wire w904;
	wire w905;
	wire w906;
	wire w907;
	wire w908;
	wire w909;
	wire w910;
	wire w911;
	wire w912;
	wire w913;
	wire w914;
	wire w915;
	wire w916;
	wire w917;
	wire w918;
	wire w919;
	wire w920;
	wire w921;
	wire w922;
	wire w923;
	wire w924;
	wire w925;
	wire w926;
	wire w927;
	wire w928;
	wire w929;
	wire w930;
	wire w931;
	wire w932;
	wire w933;
	wire w934;
	wire w935;
	wire w936;
	wire w937;
	wire w938;
	wire w939;
	wire w940;
	wire w941;
	wire w942;
	wire w943;
	wire w944;
	wire w945;
	wire w946;
	wire w947;
	wire w948;
	wire w949;
	wire w950;
	wire w951;
	wire w952;
	wire w953;
	wire w954;
	wire w955;
	wire w956;
	wire w957;
	wire w958;
	wire w959;
	wire w960;
	wire w961;
	wire w962;
	wire w963;
	wire w964;
	wire w965;
	wire w966;
	wire w967;
	wire w968;
	wire w969;
	wire w970;
	wire w971;
	wire w972;
	wire w973;

	assign n_tm_bp_cys = w760;
	assign tm_bp_cys = w211;
	assign n_sp_bp_mrd = w548;
	assign md[5] = w309;
	assign md[2] = w121;
	assign md[1] = w549;
	assign md[7] = w120;
	assign w764 = arb_fexx_ffxx;
	assign md[6] = w550;
	assign md[3] = w217;
	assign w551 = a[12];
	assign w589 = a[11];
	assign w590 = a[9];
	assign w331 = a[8];
	assign md[0] = w330;
	assign w591 = a[10];
	assign sp_bp_cys = w123;
	assign ppu_int_vbl = w378;
	assign ppu_int_stat = w377;
	assign w570 = a[4];
	assign w571 = vram_to_oam;
	assign ff46 = w637;
	assign w128 = ffxx;
	assign w129 = a[3];
	assign w912 = a[0];
	assign w130 = a[1];
	assign nma[8] = w126;
	assign w127 = a[6];
	assign ppu_mode3 = w230;
	assign w134 = a[7];
	assign nma[7] = w135;
	assign w133 = a[5];
	assign w132 = a[2];
	assign nma[1] = w131;
	assign w136 = n_ppu_hard_reset;
	assign nma[9] = w562;
	assign fexx = w817;
	assign nma[0] = w271;
	assign ff43 = w843;
	assign nma[4] = w513;
	assign nma[12] = w65;
	assign nma[6] = w270;
	assign nma[5] = w49;
	assign ff42 = w269;
	assign nma[11] = w48;
	assign w59 = ppu_rd;
	assign nma[10] = w60;
	assign w152 = ppu_wr;
	assign w153 = sprite_x_flip;
	assign w846 = n_dma_phi;
	assign n_dma_phi2_latched = w74;
	assign nma[3] = w276;
	assign nma[2] = w154;
	assign w616 = sprite_x_match;
	assign oam_mode3_bl_pch = w223;
	assign bp_sel = w222;
	assign w818 = FF43_D1;
	assign v[7] = w77;
	assign bp_cy = w209;
	assign tm_cy = w210;
	assign w11 = FF43_D0;
	assign d[4] = w68;
	assign w317 = n_ppu_clk;
	assign d[7] = w79;
	assign w821 = FF43_D2;
	assign h[3] = w171;
	assign v[6] = w172;
	assign d[1] = w12;
	assign d[3] = w52;
	assign d[6] = w248;
	assign d[2] = w91;
	assign d[0] = w13;
	assign d[5] = w339;
	assign CONST0 = w14;
	assign v[4] = w280;
	assign v[0] = w251;
	assign h[4] = w808;
	assign h[6] = w373;
	assign h[7] = w620;
	assign FF40_D3 = w54;
	assign FF40_D2 = w55;
	assign in_window = w145;
	assign h[5] = w547;
	assign w844 = h_restart;
	assign oam_mode3_nrd = w337;
	assign v[3] = w254;
	assign ppu1_ma0 = w243;
	assign v[2] = w244;
	assign h[2] = w367;
	assign oam_rd_ck = w285;
	assign v[1] = w284;
	assign v[5] = w359;
	assign oam_xattr_latch_cck = w360;
	assign FF40_D1 = w822;
	assign oam_addr_ck = w492;
	assign h[0] = w493;
	assign w366 = ppu_mode2;
	assign h[1] = w517;
	assign vbl = w953;
	assign w529 = stop_oam_eval;
	assign w198 = obj_color;
	assign vclk2 = w683;
	assign w523 = obj_prio;
	assign obj_prio_ck = w291;
	assign n_ppu_reset = w148;
	assign w365 = ppu_clk;
	assign n_ma[11] = w580;
	assign n_ma[9] = w581;
	assign n_ma[8] = w790;
	assign n_lcd_cpl = w776;
	assign n_lcd_ld1 = w4;
	assign n_lcd_cp = w5;
	assign n_lcd_st = w527;
	assign n_lcd_ld0 = w526;
	assign n_lcd_cpg = w943;
	assign n_ma[10] = w62;
	assign n_ma[12] = w63;
	assign n_lcd_fr = w418;
	assign n_lcd_s = w419;
	assign n_ma[6] = w469;
	assign n_ma[5] = w51;
	assign n_ma[7] = w510;
	assign n_ma[3] = w278;
	assign n_ma[2] = w156;
	assign n_ma[4] = w468;
	assign n_ma[1] = w387;
	assign n_ma[0] = w796;
	assign md[4] = w216;

	// Instances

	dmg_not g1 (.a(w759), .x(w323) );
	dmg_not g2 (.a(w215), .x(w918) );
	dmg_not g3 (.a(w322), .x(w324) );
	dmg_not g4 (.a(w662), .x(w661) );
	dmg_not g5 (.a(w660), .x(w659) );
	dmg_not g6 (.a(w329), .x(w328) );
	dmg_not g7 (.a(w218), .x(w119) );
	dmg_not g8 (.a(w315), .x(w756) );
	dmg_not g9 (.a(w219), .x(w218) );
	dmg_not g10 (.a(w318), .x(w166) );
	dmg_not g11 (.a(w465), .x(w466) );
	dmg_not g12 (.a(w230), .x(w663) );
	dmg_not g13 (.a(w855), .x(w95) );
	dmg_not g14 (.a(w801), .x(w93) );
	dmg_not g15 (.a(w317), .x(w596) );
	dmg_not g16 (.a(w93), .x(w92) );
	dmg_not g17 (.a(w148), .x(w406) );
	dmg_not g18 (.a(w406), .x(w421) );
	dmg_not g19 (.a(w198), .x(w940) );
	dmg_not g20 (.a(w108), .x(w728) );
	dmg_not g21 (.a(w198), .x(w769) );
	dmg_not g22 (.a(w416), .x(w933) );
	dmg_not g23 (.a(w19), .x(w434) );
	dmg_not g24 (.a(w433), .x(w187) );
	dmg_not g25 (.a(w28), .x(w27) );
	dmg_not g26 (.a(w18), .x(w932) );
	dmg_not g27 (.a(w396), .x(w345) );
	dmg_not g28 (.a(w22), .x(w21) );
	dmg_not g29 (.a(w931), .x(w390) );
	dmg_not g30 (.a(w201), .x(w200) );
	dmg_not g31 (.a(w16), .x(w441) );
	dmg_not g32 (.a(w440), .x(w17) );
	dmg_not g33 (.a(w393), .x(w392) );
	dmg_not g34 (.a(w391), .x(w394) );
	dmg_not g35 (.a(w198), .x(w524) );
	dmg_not g36 (.a(w20), .x(w483) );
	dmg_not g37 (.a(w110), .x(w111) );
	dmg_not g38 (.a(w455), .x(w454) );
	dmg_not g39 (.a(w881), .x(w880) );
	dmg_not g40 (.a(w293), .x(w410) );
	dmg_not g41 (.a(w423), .x(w744) );
	dmg_not g42 (.a(w942), .x(w624) );
	dmg_not g43 (.a(w622), .x(w623) );
	dmg_not g44 (.a(w147), .x(w146) );
	dmg_not g45 (.a(w629), .x(w802) );
	dmg_not g46 (.a(w458), .x(w457) );
	dmg_not g47 (.a(w461), .x(w459) );
	dmg_not g48 (.a(w854), .x(w221) );
	dmg_not g49 (.a(w326), .x(w325) );
	dmg_not g50 (.a(w118), .x(w313) );
	dmg_not g51 (.a(w213), .x(w212) );
	dmg_not g52 (.a(w578), .x(w548) );
	dmg_not g53 (.a(w46), .x(w45) );
	dmg_not g54 (.a(w761), .x(w960) );
	dmg_not g55 (.a(w762), .x(w853) );
	dmg_not g56 (.a(w765), .x(w552) );
	dmg_not g57 (.a(w851), .x(w910) );
	dmg_not g58 (.a(w499), .x(w500) );
	dmg_not g59 (.a(w148), .x(w531) );
	dmg_not g60 (.a(w48), .x(w579) );
	dmg_not g61 (.a(w626), .x(w628) );
	dmg_not g62 (.a(w626), .x(w627) );
	dmg_not g63 (.a(w65), .x(w64) );
	dmg_not g64 (.a(w958), .x(w959) );
	dmg_not g65 (.a(w60), .x(w61) );
	dmg_not g66 (.a(w597), .x(w598) );
	dmg_not g67 (.a(w597), .x(w609) );
	dmg_not g68 (.a(w198), .x(w944) );
	dmg_not g69 (.a(w446), .x(w34) );
	dmg_not g70 (.a(w444), .x(w936) );
	dmg_not g71 (.a(w198), .x(w786) );
	dmg_not g72 (.a(w717), .x(w199) );
	dmg_not g73 (.a(w701), .x(w697) );
	dmg_not g74 (.a(w706), .x(w699) );
	dmg_not g75 (.a(w702), .x(w698) );
	dmg_not g76 (.a(w401), .x(w789) );
	dmg_not g77 (.a(w707), .x(w672) );
	dmg_not g78 (.a(w198), .x(w945) );
	dmg_not g79 (.a(w523), .x(w712) );
	dmg_not g80 (.a(w193), .x(w194) );
	dmg_not g81 (.a(w523), .x(w687) );
	dmg_not g82 (.a(w647), .x(w450) );
	dmg_not g83 (.a(w109), .x(w108) );
	dmg_not g84 (.a(w228), .x(w861) );
	dmg_not g85 (.a(w230), .x(w594) );
	dmg_not g86 (.a(w175), .x(w206) );
	dmg_not g87 (.a(w148), .x(w644) );
	dmg_not g88 (.a(w171), .x(w375) );
	dmg_not g89 (.a(w650), .x(w376) );
	dmg_not g90 (.a(w652), .x(w653) );
	dmg_not g91 (.a(w180), .x(w181) );
	dmg_not g92 (.a(w653), .x(w654) );
	dmg_not g93 (.a(w596), .x(w164) );
	dmg_not g94 (.a(w592), .x(w906) );
	dmg_not g95 (.a(w561), .x(w962) );
	dmg_not g96 (.a(w145), .x(w794) );
	dmg_not g97 (.a(w266), .x(w265) );
	dmg_not g98 (.a(w235), .x(w162) );
	dmg_not g99 (.a(w563), .x(w264) );
	dmg_not g100 (.a(w793), .x(w263) );
	dmg_not g101 (.a(w58), .x(w57) );
	dmg_not g102 (.a(w920), .x(w67) );
	dmg_not g103 (.a(w280), .x(w967) );
	dmg_not g104 (.a(w251), .x(w966) );
	dmg_not g105 (.a(w72), .x(w71) );
	dmg_not g106 (.a(w599), .x(w835) );
	dmg_not g107 (.a(w32), .x(w823) );
	dmg_not g108 (.a(w303), .x(w302) );
	dmg_not g109 (.a(w353), .x(w351) );
	dmg_not g110 (.a(w354), .x(w352) );
	dmg_not g111 (.a(w439), .x(w353) );
	dmg_not g112 (.a(w690), .x(w691) );
	dmg_not g113 (.a(w691), .x(w448) );
	dmg_not g114 (.a(w523), .x(w826) );
	dmg_not g115 (.a(w523), .x(w949) );
	dmg_not g116 (.a(w69), .x(w70) );
	dmg_not g117 (.a(w523), .x(w834) );
	dmg_not g118 (.a(w523), .x(w832) );
	dmg_not g119 (.a(w31), .x(w30) );
	dmg_not g120 (.a(w839), .x(w69) );
	dmg_not g121 (.a(w955), .x(w341) );
	dmg_not g122 (.a(w291), .x(w36) );
	dmg_not g123 (.a(w523), .x(w682) );
	dmg_not g124 (.a(w364), .x(w363) );
	dmg_not g125 (.a(w365), .x(w364) );
	dmg_not g126 (.a(w523), .x(w684) );
	dmg_not g127 (.a(w137), .x(w82) );
	dmg_not g128 (.a(w84), .x(w83) );
	dmg_not g129 (.a(w363), .x(w362) );
	dmg_not g130 (.a(w361), .x(w360) );
	dmg_not g131 (.a(w359), .x(w358) );
	dmg_not g132 (.a(w172), .x(w335) );
	dmg_not g133 (.a(w77), .x(w78) );
	dmg_not g134 (.a(w254), .x(w336) );
	dmg_not g135 (.a(w338), .x(w337) );
	dmg_not g136 (.a(w284), .x(w283) );
	dmg_not g137 (.a(w846), .x(w150) );
	dmg_not g138 (.a(w84), .x(w85) );
	dmg_not g139 (.a(w85), .x(w535) );
	dmg_not g140 (.a(w844), .x(w537) );
	dmg_not g141 (.a(w224), .x(w223) );
	dmg_not g142 (.a(w619), .x(w618) );
	dmg_not g143 (.a(w616), .x(w617) );
	dmg_not g144 (.a(w137), .x(w138) );
	dmg_not g145 (.a(w221), .x(w222) );
	dmg_not g146 (.a(w334), .x(w273) );
	dmg_not g147 (.a(w132), .x(w793) );
	dmg_not g148 (.a(w130), .x(w563) );
	dmg_not g149 (.a(w129), .x(w235) );
	dmg_not g150 (.a(w912), .x(w266) );
	dmg_not g151 (.a(w126), .x(w791) );
	dmg_not g152 (.a(w914), .x(w370) );
	dmg_not g153 (.a(w534), .x(w88) );
	dmg_not g154 (.a(w294), .x(w293) );
	dmg_not g155 (.a(w260), .x(w259) );
	dmg_not g156 (.a(w159), .x(w158) );
	dmg_not g157 (.a(w562), .x(w582) );
	dmg_not g158 (.a(w295), .x(w110) );
	dmg_not g159 (.a(w71), .x(w247) );
	dmg_not g160 (.a(w711), .x(w708) );
	dmg_not g161 (.a(w397), .x(w700) );
	dmg_not g162 (.a(w928), .x(w398) );
	dmg_not g163 (.a(w402), .x(w788) );
	dmg_not g164 (.a(w694), .x(w354) );
	dmg_not g165 (.a(w198), .x(w787) );
	dmg_not g166 (.a(w689), .x(w690) );
	dmg_not g167 (.a(w723), .x(w722) );
	dmg_not g168 (.a(w198), .x(w860) );
	dmg_not g169 (.a(w665), .x(w859) );
	dmg_not g170 (.a(w509), .x(w968) );
	dmg_not g171 (.a(w448), .x(w307) );
	dmg_not g172 (.a(w693), .x(w305) );
	dmg_not g173 (.a(w306), .x(w946) );
	dmg_not g174 (.a(w33), .x(w865) );
	dmg_not g175 (.a(w35), .x(w304) );
	dmg_not g176 (.a(w664), .x(w455) );
	dmg_not g177 (.a(w177), .x(w652) );
	dmg_not g178 (.a(w633), .x(w383) );
	dmg_not g179 (.a(w653), .x(w498) );
	dmg_not g180 (.a(w183), .x(w165) );
	dmg_not g181 (.a(w128), .x(w847) );
	dmg_not g182 (.a(w558), .x(w584) );
	dmg_not g183 (.a(w230), .x(w8) );
	dmg_not g184 (.a(w506), .x(w507) );
	dmg_not g185 (.a(w148), .x(w176) );
	dmg_not g186 (.a(w609), .x(w608) );
	dmg_not g187 (.a(w610), .x(w528) );
	dmg_not g188 (.a(w738), .x(w736) );
	dmg_not g189 (.a(w735), .x(w175) );
	dmg_not g190 (.a(w202), .x(w881) );
	dmg_not g191 (.a(w880), .x(w446) );
	dmg_not g192 (.a(w694), .x(w393) );
	dmg_not g193 (.a(w439), .x(w391) );
	dmg_not g194 (.a(w435), .x(w104) );
	dmg_not g195 (.a(w244), .x(w258) );
	dmg_not g196 (.a(w276), .x(w277) );
	dmg_not g197 (.a(w154), .x(w155) );
	dmg_not g198 (.a(w88), .x(w811) );
	dmg_not g199 (.a(w270), .x(w888) );
	dmg_not g200 (.a(w49), .x(w50) );
	dmg_not g201 (.a(w317), .x(w812) );
	dmg_not g202 (.a(w317), .x(w890) );
	dmg_not g203 (.a(w317), .x(w655) );
	dmg_not g204 (.a(w271), .x(w795) );
	dmg_not g205 (.a(w513), .x(w514) );
	dmg_not g206 (.a(w135), .x(w511) );
	dmg_not g207 (.a(w131), .x(w386) );
	dmg_not g208 (.a(w220), .x(w219) );
	dmg_not g209 (.a(w759), .x(w760) );
	dmg_dffsr g210 (.nset1(w799), .nset2(w799), .clk(w44), .nres(w930), .d(w25), .q(w716) );
	dmg_dffsr g211 (.nset1(w24), .nset2(w24), .clk(w44), .nres(w395), .d(w23), .q(w25) );
	dmg_dffsr g212 (.nset1(w29), .nset2(w29), .clk(w44), .nres(w970), .d(w470), .q(w28) );
	dmg_dffsr g213 (.nset1(w214), .nset2(w214), .clk(w44), .nres(w114), .d(w320), .q(w115) );
	dmg_dffsr g214 (.nset1(w117), .nset2(w117), .clk(w44), .nres(w753), .d(w116), .q(w752) );
	dmg_dffsr g215 (.nset1(w754), .nset2(w754), .clk(w44), .nres(w814), .d(w916), .q(w917) );
	dmg_dffsr g216 (.nset1(w195), .nset2(w195), .clk(w44), .nres(w772), .d(w196), .q(w771) );
	dmg_dffsr g217 (.nset1(w15), .nset2(w15), .clk(w44), .nres(w934), .d(w14), .q(w778) );
	dmg_dffsr g218 (.nset1(w935), .nset2(w935), .clk(w44), .nres(w782), .d(w14), .q(w779) );
	dmg_dffsr g219 (.nset1(w720), .nset2(w720), .clk(w44), .nres(w719), .d(w442), .q(w37) );
	dmg_dffsr g220 (.nset1(w670), .nset2(w670), .clk(w44), .nres(w784), .d(w669), .q(w724) );
	dmg_dffsr g221 (.nset1(w938), .nset2(w938), .clk(w44), .nres(w667), .d(w14), .q(w668) );
	dmg_dffsr g222 (.nset1(w586), .nset2(w586), .clk(w44), .nres(w763), .d(w585), .q(w852) );
	dmg_dffsr g223 (.nset1(w555), .nset2(w555), .clk(w44), .nres(w911), .d(w554), .q(w556) );
	dmg_dffsr g224 (.nset1(w903), .nset2(w903), .clk(w44), .nres(w904), .d(w902), .q(w559) );
	dmg_dffsr g225 (.nset1(w907), .nset2(w907), .clk(w44), .nres(w901), .d(w14), .q(w902) );
	dmg_dffsr g226 (.nset1(w676), .nset2(w676), .clk(w44), .nres(w677), .d(w675), .q(w678) );
	dmg_dffsr g227 (.nset1(w715), .nset2(w715), .clk(w44), .nres(w833), .d(w716), .q(w190) );
	dmg_dffsr g228 (.nset1(w921), .nset2(w921), .clk(w44), .nres(w927), .d(w189), .q(w923) );
	dmg_dffsr g229 (.nset1(w191), .nset2(w191), .clk(w44), .nres(w922), .d(w190), .q(w192) );
	dmg_dffsr g230 (.nset1(w837), .nset2(w837), .clk(w44), .nres(w838), .d(w39), .q(w40) );
	dmg_dffsr g231 (.nset1(w474), .nset2(w474), .clk(w44), .nres(w836), .d(w473), .q(w43) );
	dmg_dffsr g232 (.nset1(w301), .nset2(w301), .clk(w44), .nres(w681), .d(w680), .q(w300) );
	dmg_dffsr g233 (.nset1(w679), .nset2(w679), .clk(w44), .nres(w952), .d(w678), .q(w680) );
	dmg_dffsr g234 (.nset1(w673), .nset2(w673), .clk(w44), .nres(w710), .d(w38), .q(w39) );
	dmg_dffsr g235 (.nset1(w924), .nset2(w924), .clk(w44), .nres(w713), .d(w923), .q(w675) );
	dmg_dffsr g236 (.nset1(w948), .nset2(w948), .clk(w44), .nres(w472), .d(w192), .q(w473) );
	dmg_dffsr g237 (.nset1(w688), .nset2(w688), .clk(w44), .nres(w947), .d(w40), .q(w41) );
	dmg_dffsr g238 (.nset1(w863), .nset2(w863), .clk(w44), .nres(w864), .d(w41), .q(w42) );
	dmg_dffsr g239 (.nset1(w186), .nset2(w186), .clk(w44), .nres(w188), .d(w47), .q(w189) );
	dmg_dffsr g240 (.nset1(w299), .nset2(w299), .clk(w44), .nres(w686), .d(w300), .q(w298) );
	dmg_dffsr g241 (.nset1(w297), .nset2(w297), .clk(w44), .nres(w685), .d(w298), .q(w296) );
	dmg_dffsr g242 (.nset1(w577), .nset2(w577), .clk(w44), .nres(w553), .d(w588), .q(w554) );
	dmg_dffsr g243 (.nset1(w560), .nset2(w560), .clk(w44), .nres(w961), .d(w559), .q(w585) );
	dmg_dffsr g244 (.nset1(w557), .nset2(w557), .clk(w44), .nres(w141), .d(w556), .q(w140) );
	dmg_dffsr g245 (.nset1(w587), .nset2(w587), .clk(w44), .nres(w905), .d(w852), .q(w588) );
	dmg_dffsr g246 (.nset1(w705), .nset2(w705), .clk(w44), .nres(w704), .d(w668), .q(w669) );
	dmg_dffsr g247 (.nset1(w725), .nset2(w725), .clk(w44), .nres(w726), .d(w724), .q(w785) );
	dmg_dffsr g248 (.nset1(w721), .nset2(w721), .clk(w44), .nres(w718), .d(w37), .q(w38) );
	dmg_dffsr g249 (.nset1(w671), .nset2(w671), .clk(w44), .nres(w197), .d(w785), .q(w196) );
	dmg_dffsr g250 (.nset1(w777), .nset2(w777), .clk(w44), .nres(w443), .d(w778), .q(w442) );
	dmg_dffsr g251 (.nset1(w310), .nset2(w310), .clk(w44), .nres(w112), .d(w752), .q(w751) );
	dmg_dffsr g252 (.nset1(w321), .nset2(w321), .clk(w44), .nres(w757), .d(w319), .q(w320) );
	dmg_dffsr g253 (.nset1(w658), .nset2(w658), .clk(w44), .nres(w657), .d(w115), .q(w116) );
	dmg_dffsr g254 (.nset1(w314), .nset2(w314), .clk(w44), .nres(w755), .d(w917), .q(w319) );
	dmg_dffsr g255 (.nset1(w327), .nset2(w327), .clk(w44), .nres(w758), .d(w14), .q(w916) );
	dmg_dffsr g256 (.nset1(w471), .nset2(w471), .clk(w44), .nres(w770), .d(w771), .q(w470) );
	dmg_dffsr g257 (.nset1(w780), .nset2(w780), .clk(w44), .nres(w783), .d(w779), .q(w23) );
	dmg_dffr g258 (.clk(w655), .nr1(w143), .nr2(w143), .d(w166), .nq(w316) );
	dmg_dffr g259 (.clk(w464), .nr1(w143), .nr2(w143), .d(w463), .nq(w463), .q(w465) );
	dmg_dffr g260 (.clk(w317), .nr1(w230), .nr2(w230), .d(w465), .q(w467) );
	dmg_dffr g261 (.clk(w409), .nr1(w256), .nr2(w256), .d(w257), .nq(w257), .q(w244) );
	dmg_dffr g262 (.clk(w257), .nr1(w256), .nr2(w256), .d(w255), .nq(w255), .q(w254) );
	dmg_dffr g263 (.clk(w255), .nr1(w256), .nr2(w256), .d(w279), .nq(w279), .q(w280) );
	dmg_dffr g264 (.clk(w279), .nr1(w256), .nr2(w256), .d(w408), .nq(w408), .q(w359) );
	dmg_dffr g265 (.clk(w489), .nr1(w256), .nr2(w256), .d(w76), .nq(w76), .q(w77) );
	dmg_dffr g266 (.clk(w692), .nr1(w421), .nr2(w421), .d(w969), .nq(w969) );
	dmg_dffr g267 (.clk(w933), .nr1(w421), .nr2(w421), .d(w692), .nq(w692) );
	dmg_dffr g268 (.clk(w734), .nr1(w421), .nr2(w421), .d(w733), .nq(w733), .q(w956) );
	dmg_dffr g269 (.clk(w509), .nr1(w421), .nr2(w421), .d(w416), .nq(w173), .q(w174) );
	dmg_dffr g270 (.clk(w317), .nr1(w148), .nr2(w148), .d(w147), .nq(w630) );
	dmg_dffr g271 (.clk(w812), .nr1(w230), .nr2(w230), .d(w804), .nq(w803) );
	dmg_dffr g272 (.clk(w890), .nr1(w148), .nr2(w148), .d(w168), .q(w532) );
	dmg_dffr g273 (.clk(w317), .nr1(w167), .nr2(w167), .d(w166), .q(w868) );
	dmg_dffr g274 (.clk(w462), .nr1(w143), .nr2(w143), .d(w915), .nq(w915), .q(w854) );
	dmg_dffr g275 (.clk(w317), .nr1(w230), .nr2(w230), .d(w750), .q(w900) );
	dmg_dffr g276 (.clk(w626), .nr1(w230), .nr2(w230), .d(w625), .nq(w909), .q(w750) );
	dmg_dffr g277 (.clk(w878), .nr1(w501), .nr2(w501), .d(w895), .nq(w895), .q(w876) );
	dmg_dffr g278 (.clk(w505), .nr1(w501), .nr2(w501), .d(w878), .nq(w878), .q(w877) );
	dmg_dffr g279 (.clk(w502), .nr1(w501), .nr2(w501), .d(w505), .nq(w505), .q(w504) );
	dmg_dffr g280 (.clk(w509), .nr1(w246), .nr2(w246), .d(w736), .q(w546) );
	dmg_dffr g281 (.clk(w968), .nr1(w421), .nr2(w421), .d(w727), .q(w416) );
	dmg_dffr g282 (.clk(w404), .nr1(w405), .nr2(w405), .d(w703), .nq(w703), .q(w928) );
	dmg_dffr g283 (.clk(w926), .nr1(w405), .nr2(w405), .d(w674), .nq(w674), .q(w702) );
	dmg_dffr g284 (.clk(w674), .nr1(w405), .nr2(w405), .d(w714), .nq(w714), .q(w706) );
	dmg_dffr g285 (.clk(w925), .nr1(w405), .nr2(w405), .d(w403), .nq(w403), .q(w402) );
	dmg_dffr g286 (.clk(w596), .nr1(w47), .nr2(w47), .d(w228), .nq(w239), .q(w204) );
	dmg_dffr g287 (.clk(w815), .nr1(w816), .nr2(w816), .d(w227), .nq(w227), .q(w228) );
	dmg_dffr g288 (.clk(w227), .nr1(w816), .nr2(w816), .d(w964), .nq(w964), .q(w522) );
	dmg_dffr g289 (.clk(w964), .nr1(w816), .nr2(w816), .d(w965), .nq(w965), .q(w226) );
	dmg_dffr g290 (.clk(w375), .nr1(w495), .nr2(w495), .d(w894), .q(w547) );
	dmg_dffr g291 (.clk(w375), .nr1(w495), .nr2(w495), .d(w871), .q(w373) );
	dmg_dffr g292 (.clk(w375), .nr1(w495), .nr2(w495), .d(w874), .nq(w874), .q(w808) );
	dmg_dffr g293 (.clk(w164), .nr1(w230), .nr2(w230), .d(w522), .q(w521) );
	dmg_dffr g294 (.clk(w634), .nr1(w383), .nr2(w383), .d(w639), .nq(w639), .q(w640) );
	dmg_dffr g295 (.clk(w639), .nr1(w383), .nr2(w383), .d(w384), .nq(w384), .q(w963) );
	dmg_dffr g296 (.clk(w384), .nr1(w383), .nr2(w383), .d(w575), .nq(w575), .q(w576) );
	dmg_dffr g297 (.clk(w575), .nr1(w383), .nr2(w383), .d(w124), .nq(w124), .q(w125) );
	dmg_dffr g298 (.clk(w124), .nr1(w383), .nr2(w383), .d(w574), .nq(w574), .q(w573) );
	dmg_dffr g299 (.clk(w379), .nr1(w273), .nr2(w273), .d(w274), .nq(w274), .q(w275) );
	dmg_dffr g300 (.clk(w566), .nr1(w273), .nr2(w273), .d(w379), .nq(w379), .q(w380) );
	dmg_dffr g301 (.clk(w564), .nr1(w273), .nr2(w273), .d(w566), .nq(w566), .q(w565) );
	dmg_dffr g302 (.clk(w583), .nr1(w273), .nr2(w273), .d(w564), .nq(w564), .q(w272) );
	dmg_dffr g303 (.clk(w363), .nr1(w148), .nr2(w148), .d(w288), .nq(w288) );
	dmg_dffr g304 (.clk(w362), .nr1(w148), .nr2(w148), .d(w288), .nq(w287), .q(w286) );
	dmg_dffr g305 (.clk(w150), .nr1(w138), .nr2(w138), .d(w149) );
	dmg_dffr g306 (.clk(w44), .nr1(w495), .nr2(w495), .d(w825), .q(w367) );
	dmg_dffr g307 (.clk(w44), .nr1(w495), .nr2(w495), .d(w518), .q(w171) );
	dmg_dffr g308 (.clk(w44), .nr1(w495), .nr2(w495), .d(w494), .nq(w494), .q(w493) );
	dmg_dffr g309 (.clk(w274), .nr1(w273), .nr2(w273), .d(w636), .nq(w636), .q(w635) );
	dmg_dffr g310 (.clk(w794), .nr1(w383), .nr2(w383), .d(w638), .nq(w638), .q(w385) );
	dmg_dffr g311 (.clk(w638), .nr1(w383), .nr2(w383), .d(w382), .nq(w382), .q(w381) );
	dmg_dffr g312 (.clk(w382), .nr1(w383), .nr2(w383), .d(w634), .nq(w634), .q(w332) );
	dmg_dffr g313 (.clk(w317), .nr1(w495), .nr2(w495), .d(w496), .q(w615) );
	dmg_dffr g314 (.clk(w164), .nr1(w230), .nr2(w230), .d(w521), .nq(w242), .q(w241) );
	dmg_dffr g315 (.clk(w288), .nr1(w148), .nr2(w148), .d(w862), .nq(w862) );
	dmg_dffr g316 (.clk(w403), .nr1(w405), .nr2(w405), .d(w404), .nq(w404), .q(w397) );
	dmg_dffr g317 (.clk(w703), .nr1(w405), .nr2(w405), .d(w926), .nq(w926), .q(w701) );
	dmg_dffr g318 (.clk(w968), .nr1(w421), .nr2(w421), .d(w929), .q(w666) );
	dmg_dffr g319 (.clk(w509), .nr1(w405), .nr2(w405), .d(w925), .nq(w925), .q(w401) );
	dmg_dffr g320 (.clk(w509), .nr1(w148), .nr2(w148), .d(w959), .q(w749) );
	dmg_dffr g321 (.clk(w44), .nr1(w495), .nr2(w495), .d(w971), .q(w517) );
	dmg_dffr g322 (.clk(w596), .nr1(w230), .nr2(w230), .d(w241), .q(w229) );
	dmg_dffr g323 (.clk(w375), .nr1(w495), .nr2(w495), .d(w892), .q(w620) );
	dmg_dffr g324 (.clk(w317), .nr1(w148), .nr2(w148), .d(w177), .q(w875) );
	dmg_dffr g325 (.clk(w164), .nr1(w47), .nr2(w47), .d(w869), .q(w185) );
	dmg_dffr g326 (.clk(w596), .nr1(w47), .nr2(w47), .d(w185), .nq(w184) );
	dmg_dffr g327 (.clk(w655), .nr1(w167), .nr2(w167), .d(w868), .q(w179) );
	dmg_dffr g328 (.clk(w317), .nr1(w230), .nr2(w230), .d(w179), .q(w867) );
	dmg_dffr g329 (.clk(w628), .nr1(w230), .nr2(w230), .d(w507), .q(w804) );
	dmg_dffr g330 (.clk(w627), .nr1(w148), .nr2(w148), .d(w624), .q(w168) );
	dmg_dffr g331 (.clk(w628), .nr1(w230), .nr2(w230), .d(w171), .q(w426) );
	dmg_dffr g332 (.clk(w174), .nr1(w421), .nr2(w421), .d(w953), .nq(w735), .q(w734) );
	dmg_dffr g333 (.clk(w173), .nr1(w421), .nr2(w421), .d(w540), .q(w407) );
	dmg_dffr g334 (.clk(w173), .nr1(w421), .nr2(w421), .d(w422), .q(w420) );
	dmg_dffr g335 (.clk(w408), .nr1(w256), .nr2(w256), .d(w489), .nq(w489), .q(w172) );
	dmg_dffr g336 (.clk(w416), .nr1(w256), .nr2(w256), .d(w252), .nq(w252), .q(w251) );
	dmg_dffr g337 (.clk(w252), .nr1(w256), .nr2(w256), .d(w409), .nq(w409), .q(w284) );
	dmg_dffr g338 (.clk(w463), .nr1(w143), .nr2(w143), .d(w462), .nq(w462), .q(w461) );
	dmg_nand g339 (.a(w113), .b(w322), .x(w321) );
	dmg_nand g340 (.a(w324), .b(w113), .x(w757) );
	dmg_nand g341 (.a(w113), .b(w660), .x(w658) );
	dmg_nand g342 (.a(w659), .b(w113), .x(w657) );
	dmg_nand g343 (.a(w113), .b(w329), .x(w327) );
	dmg_nand g344 (.a(w328), .b(w113), .x(w758) );
	dmg_nand g345 (.a(w756), .b(w113), .x(w755) );
	dmg_nand g346 (.a(w113), .b(w315), .x(w314) );
	dmg_nand g347 (.a(w317), .b(w318), .x(w464) );
	dmg_nand g348 (.a(w198), .b(w30), .x(w29) );
	dmg_nand g349 (.a(w940), .b(w30), .x(w970) );
	dmg_nand g350 (.a(w198), .b(w305), .x(w471) );
	dmg_nand g351 (.a(w769), .b(w305), .x(w770) );
	dmg_nand g352 (.a(w28), .b(w435), .x(w931) );
	dmg_nand g353 (.a(w18), .b(w17), .x(w24) );
	dmg_nand g354 (.a(w932), .b(w17), .x(w395) );
	dmg_nand g355 (.a(w27), .b(w435), .x(w396) );
	dmg_nand g356 (.a(w200), .b(w199), .x(w930) );
	dmg_nand g357 (.a(w459), .b(w221), .x(w458) );
	dmg_nand g358 (.a(w113), .b(w326), .x(w754) );
	dmg_nand g359 (.a(w325), .b(w113), .x(w814) );
	dmg_nand g360 (.a(w113), .b(w118), .x(w117) );
	dmg_nand g361 (.a(w313), .b(w113), .x(w753) );
	dmg_nand g362 (.a(w113), .b(w213), .x(w310) );
	dmg_nand g363 (.a(w212), .b(w113), .x(w112) );
	dmg_nand g364 (.a(w142), .b(w46), .x(w577) );
	dmg_nand g365 (.a(w142), .b(w561), .x(w560) );
	dmg_nand g366 (.a(w142), .b(w761), .x(w555) );
	dmg_nand g367 (.a(w584), .b(w142), .x(w141) );
	dmg_nand g368 (.a(w142), .b(w558), .x(w557) );
	dmg_nand g369 (.a(w142), .b(w765), .x(w586) );
	dmg_nand g370 (.a(w142), .b(w851), .x(w587) );
	dmg_nand g371 (.a(w847), .b(w764), .x(w848) );
	dmg_nand g372 (.a(w972), .b(w739), .x(w738) );
	dmg_nand g373 (.a(w665), .b(w21), .x(w777) );
	dmg_nand g374 (.a(w859), .b(w21), .x(w443) );
	dmg_nand g375 (.a(w786), .b(w672), .x(w197) );
	dmg_nand g376 (.a(w198), .b(w672), .x(w671) );
	dmg_nand g377 (.a(w723), .b(w199), .x(w721) );
	dmg_nand g378 (.a(w722), .b(w199), .x(w718) );
	dmg_nand g379 (.a(w787), .b(w199), .x(w726) );
	dmg_nand g380 (.a(w945), .b(w21), .x(w704) );
	dmg_nand g381 (.a(w711), .b(w672), .x(w673) );
	dmg_nand g382 (.a(w712), .b(w17), .x(w713) );
	dmg_nand g383 (.a(w523), .b(w17), .x(w924) );
	dmg_nand g384 (.a(w946), .b(w305), .x(w472) );
	dmg_nand g385 (.a(w306), .b(w305), .x(w948) );
	dmg_nand g386 (.a(w687), .b(w305), .x(w686) );
	dmg_nand g387 (.a(w33), .b(w305), .x(w688) );
	dmg_nand g388 (.a(w865), .b(w305), .x(w947) );
	dmg_nand g389 (.a(w304), .b(w30), .x(w864) );
	dmg_nand g390 (.a(w35), .b(w30), .x(w863) );
	dmg_nand g391 (.a(w523), .b(w305), .x(w299) );
	dmg_nand g392 (.a(w523), .b(w30), .x(w297) );
	dmg_nand g393 (.a(w523), .b(w187), .x(w186) );
	dmg_nand g394 (.a(w861), .b(w204), .x(w205) );
	dmg_nand g395 (.a(w226), .b(w228), .x(w595) );
	dmg_nand g396 (.a(w875), .b(w652), .x(w497) );
	dmg_nand g397 (.a(w684), .b(w30), .x(w685) );
	dmg_nand g398 (.a(w682), .b(w187), .x(w188) );
	dmg_nand g399 (.a(w834), .b(w194), .x(w681) );
	dmg_nand g400 (.a(w832), .b(w21), .x(w927) );
	dmg_nand g401 (.a(w708), .b(w672), .x(w710) );
	dmg_nand g402 (.a(w949), .b(w672), .x(w952) );
	dmg_nand g403 (.a(w826), .b(w199), .x(w677) );
	dmg_nand g404 (.a(w523), .b(w199), .x(w676) );
	dmg_nand g405 (.a(w523), .b(w672), .x(w679) );
	dmg_nand g406 (.a(w523), .b(w21), .x(w921) );
	dmg_nand g407 (.a(w709), .b(w672), .x(w833) );
	dmg_nand g408 (.a(w302), .b(w194), .x(w922) );
	dmg_nand g409 (.a(w823), .b(w194), .x(w838) );
	dmg_nand g410 (.a(w835), .b(w30), .x(w836) );
	dmg_nand g411 (.a(w523), .b(w194), .x(w301) );
	dmg_nand g412 (.a(w81), .b(w82), .x(w954) );
	dmg_nand g413 (.a(w209), .b(w145), .x(w333) );
	dmg_nand g414 (.a(w599), .b(w30), .x(w474) );
	dmg_nand g415 (.a(w32), .b(w194), .x(w837) );
	dmg_nand g416 (.a(w303), .b(w194), .x(w191) );
	dmg_nand g417 (.a(w484), .b(w672), .x(w715) );
	dmg_nand g418 (.a(w198), .b(w199), .x(w725) );
	dmg_nand g419 (.a(w198), .b(w21), .x(w705) );
	dmg_nand g420 (.a(w860), .b(w187), .x(w667) );
	dmg_nand g421 (.a(w596), .b(w595), .x(w815) );
	dmg_nand g422 (.a(w910), .b(w142), .x(w905) );
	dmg_nand g423 (.a(w906), .b(w142), .x(w901) );
	dmg_nand g424 (.a(w552), .b(w142), .x(w763) );
	dmg_nand g425 (.a(w142), .b(w762), .x(w903) );
	dmg_nand g426 (.a(w853), .b(w142), .x(w904) );
	dmg_nand g427 (.a(w960), .b(w142), .x(w911) );
	dmg_nand g428 (.a(w962), .b(w142), .x(w961) );
	dmg_nand g429 (.a(w45), .b(w142), .x(w553) );
	dmg_nand g430 (.a(w628), .b(w503), .x(w502) );
	dmg_nand g431 (.a(w198), .b(w187), .x(w938) );
	dmg_nand g432 (.a(w444), .b(w187), .x(w935) );
	dmg_nand g433 (.a(w198), .b(w17), .x(w670) );
	dmg_nand g434 (.a(w524), .b(w17), .x(w784) );
	dmg_nand g435 (.a(w441), .b(w17), .x(w719) );
	dmg_nand g436 (.a(w16), .b(w17), .x(w720) );
	dmg_nand g437 (.a(w201), .b(w199), .x(w799) );
	dmg_nand g438 (.a(w483), .b(w21), .x(w783) );
	dmg_nand g439 (.a(w20), .b(w21), .x(w780) );
	dmg_nand g440 (.a(w434), .b(w187), .x(w934) );
	dmg_nand g441 (.a(w19), .b(w187), .x(w15) );
	dmg_nand g442 (.a(w198), .b(w194), .x(w195) );
	dmg_nand g443 (.a(w918), .b(w113), .x(w114) );
	dmg_nand g444 (.a(w113), .b(w215), .x(w214) );
	dmg_latch_comp g445 (.n_ena(w218), .d(w217), .ena(w119), .q(w322) );
	dmg_latch_comp g446 (.n_ena(w218), .d(w330), .ena(w119), .q(w329) );
	dmg_latch_comp g447 (.n_ena(w218), .d(w549), .ena(w119), .q(w326) );
	dmg_latch_comp g448 (.n_ena(w218), .d(w550), .ena(w119), .q(w118) );
	dmg_latch_comp g449 (.n_ena(w218), .d(w120), .ena(w119), .q(w213) );
	dmg_latch_comp g450 (.n_ena(w446), .d(w308), .ena(w34), .q(w35) );
	dmg_latch_comp g451 (.n_ena(w446), .d(w447), .ena(w34), .q(w33) );
	dmg_latch_comp g452 (.n_ena(w446), .d(w445), .ena(w34), .q(w723) );
	dmg_latch_comp g453 (.n_ena(w448), .d(w879), .ena(w307), .q(w444) );
	dmg_latch_comp g454 (.n_ena(w446), .d(w766), .ena(w34), .q(w665) );
	dmg_latch_comp g455 (.n_ena(w448), .d(w485), .ena(w307), .q(w484) );
	dmg_latch_comp g456 (.n_ena(w446), .d(w485), .ena(w34), .q(w711) );
	dmg_latch_comp g457 (.n_ena(w448), .d(w447), .ena(w307), .q(w306) );
	dmg_latch_comp g458 (.n_ena(w446), .d(w866), .ena(w34), .q(w32) );
	dmg_latch_comp g459 (.n_ena(w448), .d(w866), .ena(w307), .q(w303) );
	dmg_latch_comp g460 (.n_ena(w448), .d(w308), .ena(w307), .q(w599) );
	dmg_latch_comp g461 (.n_ena(w448), .d(w445), .ena(w307), .q(w201) );
	dmg_latch_comp g462 (.n_ena(w446), .d(w879), .ena(w34), .q(w19) );
	dmg_latch_comp g463 (.n_ena(w448), .d(w766), .ena(w307), .q(w20) );
	dmg_latch_comp g464 (.n_ena(w448), .d(w456), .ena(w307), .q(w18) );
	dmg_latch_comp g465 (.n_ena(w446), .d(w456), .ena(w34), .q(w16) );
	dmg_latch_comp g466 (.n_ena(w218), .d(w121), .ena(w119), .q(w315) );
	dmg_latch_comp g467 (.n_ena(w218), .d(w216), .ena(w119), .q(w215) );
	dmg_latch_comp g468 (.n_ena(w218), .d(w309), .ena(w119), .q(w660) );
	dmg_not2 g469 (.a(w323), .x(w211) );
	dmg_not2 g470 (.a(w661), .x(w312) );
	dmg_not2 g471 (.a(w312), .x(w311) );
	dmg_not2 g472 (.a(w143), .x(w142) );
	dmg_not2 g473 (.a(w143), .x(w113) );
	dmg_not2 g474 (.a(w386), .x(w387) );
	dmg_not2 g475 (.a(w514), .x(w468) );
	dmg_not2 g476 (.a(w511), .x(w510) );
	dmg_not2 g477 (.a(w795), .x(w796) );
	dmg_not2 g478 (.a(w50), .x(w51) );
	dmg_not2 g479 (.a(w888), .x(w469) );
	dmg_not2 g480 (.a(w155), .x(w156) );
	dmg_not2 g481 (.a(w277), .x(w278) );
	dmg_not2 g482 (.a(w61), .x(w62) );
	dmg_not2 g483 (.a(w3), .x(w4) );
	dmg_not2 g484 (.a(w525), .x(w526) );
	dmg_not2 g485 (.a(w582), .x(w581) );
	dmg_not2 g486 (.a(w791), .x(w790) );
	dmg_not2 g487 (.a(w163), .x(w870) );
	dmg_nand g488 (.a(w142), .x(w907), .b(w592) );
	dmg_not2 g489 (.a(w593), .x(w123) );
	dmg_not2 g490 (.a(w512), .x(w572) );
	dmg_not2 g491 (.a(w568), .x(w267) );
	dmg_not2 g492 (.a(w645), .x(w646) );
	dmg_not2 g493 (.a(w137), .x(w249) );
	dmg_not2 g494 (.a(w290), .x(w291) );
	dmg_not2 g495 (.a(w137), .x(w246) );
	dmg_not2 g496 (.a(w841), .x(w840) );
	dmg_not2 g497 (.a(w954), .x(w148) );
	dmg_not2 g498 (.a(w286), .x(w285) );
	dmg_not2 g499 (.a(w288), .x(w492) );
	dmg_not2 g500 (.a(w75), .x(w74) );
	dmg_not2 g501 (.a(w242), .x(w243) );
	dmg_not2 g502 (.a(w913), .x(w73) );
	dmg_not2 g503 (.a(w842), .x(w843) );
	dmg_not2 g504 (.a(w262), .x(w261) );
	dmg_not2 g505 (.a(w268), .x(w269) );
	dmg_not2 g506 (.a(w136), .x(w137) );
	dmg_not2 g507 (.a(w237), .x(w236) );
	dmg_not2 g508 (.a(w567), .x(w637) );
	dmg_not2 g509 (.a(w161), .x(w160) );
	dmg_not2 g510 (.a(w792), .x(w533) );
	dmg_not2 g511 (.a(w234), .x(w233) );
	dmg_not2 g512 (.a(w919), .x(w292) );
	dmg_not2 g513 (.a(w776), .x(w683) );
	dmg_not2 g514 (.a(w848), .x(w817) );
	dmg_not2 g515 (.a(w497), .x(w898) );
	dmg_not2 g516 (.a(w146), .x(w145) );
	dmg_not2 g517 (.a(w858), .x(w943) );
	dmg_not2 g518 (.a(w64), .x(w63) );
	dmg_not2 g519 (.a(w579), .x(w580) );
	dmg_not2 g520 (.a(w802), .x(w891) );
	dmg_notif0 g521 (.n_ena(w95), .a(w431), .x(w339) );
	dmg_notif0 g522 (.n_ena(w95), .a(w856), .x(w13) );
	dmg_notif0 g523 (.n_ena(w95), .a(w96), .x(w91) );
	dmg_notif0 g524 (.n_ena(w95), .a(w797), .x(w79) );
	dmg_notif0 g525 (.n_ena(w95), .a(w889), .x(w248) );
	dmg_notif0 g526 (.n_ena(w95), .a(w100), .x(w52) );
	dmg_notif0 g527 (.n_ena(w95), .a(w94), .x(w68) );
	dmg_notif0 g528 (.n_ena(w95), .a(w883), .x(w12) );
	dmg_notif0 g529 (.n_ena(w370), .a(w515), .x(w13) );
	dmg_notif0 g530 (.n_ena(w370), .a(w885), .x(w52) );
	dmg_notif0 g531 (.n_ena(w259), .a(w258), .x(w91) );
	dmg_notif0 g532 (.n_ena(w158), .a(w157), .x(w52) );
	dmg_notif0 g533 (.n_ena(w450), .a(w101), .x(w52) );
	dmg_notif0 g534 (.n_ena(w450), .a(w729), .x(w68) );
	dmg_notif0 g535 (.n_ena(w450), .a(w730), .x(w79) );
	dmg_notif0 g536 (.n_ena(w450), .a(w488), .x(w339) );
	dmg_notif0 g537 (.n_ena(w450), .a(w480), .x(w248) );
	dmg_notif0 g538 (.n_ena(w236), .a(w589), .x(w48) );
	dmg_notif0 g539 (.n_ena(w236), .a(w590), .x(w562) );
	dmg_notif0 g540 (.n_ena(w236), .a(w331), .x(w126) );
	dmg_notif0 g541 (.n_ena(w236), .a(w591), .x(w60) );
	dmg_notif0 g542 (.n_ena(w236), .a(w551), .x(w65) );
	dmg_notif0 g543 (.n_ena(w67), .a(w747), .x(w91) );
	dmg_notif0 g544 (.n_ena(w67), .a(w746), .x(w13) );
	dmg_notif0 g545 (.n_ena(w67), .a(w602), .x(w52) );
	dmg_notif0 g546 (.n_ena(w67), .a(w601), .x(w68) );
	dmg_notif0 g547 (.n_ena(w450), .a(w107), .x(w13) );
	dmg_notif0 g548 (.n_ena(w450), .a(w449), .x(w91) );
	dmg_notif0 g549 (.n_ena(w333), .a(w381), .x(w154) );
	dmg_notif0 g550 (.n_ena(w333), .a(w385), .x(w131) );
	dmg_notif0 g551 (.n_ena(w333), .a(w332), .x(w276) );
	dmg_notif0 g552 (.n_ena(w572), .a(w635), .x(w513) );
	dmg_notif0 g553 (.n_ena(w57), .a(w86), .x(w13) );
	dmg_notif0 g554 (.n_ena(w57), .a(w53), .x(w52) );
	dmg_notif0 g555 (.n_ena(w57), .a(w56), .x(w91) );
	dmg_notif0 g556 (.n_ena(w259), .a(w335), .x(w248) );
	dmg_notif0 g557 (.n_ena(w259), .a(w78), .x(w79) );
	dmg_notif0 g558 (.n_ena(w259), .a(w336), .x(w52) );
	dmg_notif0 g559 (.n_ena(w259), .a(w358), .x(w339) );
	dmg_notif0 g560 (.n_ena(w259), .a(w283), .x(w12) );
	dmg_notif0 g561 (.n_ena(w341), .a(w342), .x(w13) );
	dmg_notif0 g562 (.n_ena(w341), .a(w951), .x(w91) );
	dmg_notif0 g563 (.n_ena(w341), .a(w357), .x(w52) );
	dmg_notif0 g564 (.n_ena(w341), .a(w348), .x(w79) );
	dmg_notif0 g565 (.n_ena(w341), .a(w340), .x(w339) );
	dmg_notif0 g566 (.n_ena(w341), .a(w824), .x(w248) );
	dmg_notif0 g567 (.n_ena(w341), .a(w829), .x(w68) );
	dmg_notif0 g568 (.n_ena(w341), .a(w828), .x(w12) );
	dmg_notif0 g569 (.n_ena(w57), .a(w973), .x(w12) );
	dmg_notif0 g570 (.n_ena(w57), .a(w80), .x(w79) );
	dmg_notif0 g571 (.n_ena(w236), .a(w133), .x(w49) );
	dmg_notif0 g572 (.n_ena(w236), .a(w132), .x(w154) );
	dmg_notif0 g573 (.n_ena(w236), .a(w570), .x(w513) );
	dmg_notif0 g574 (.n_ena(w236), .a(w134), .x(w135) );
	dmg_notif0 g575 (.n_ena(w236), .a(w127), .x(w270) );
	dmg_notif0 g576 (.n_ena(w333), .a(w222), .x(w271) );
	dmg_notif0 g577 (.n_ena(w236), .a(w912), .x(w271) );
	dmg_notif0 g578 (.n_ena(w236), .a(w130), .x(w131) );
	dmg_notif0 g579 (.n_ena(w572), .a(w272), .x(w271) );
	dmg_notif0 g580 (.n_ena(w236), .a(w129), .x(w276) );
	dmg_notif0 g581 (.n_ena(w572), .a(w565), .x(w131) );
	dmg_notif0 g582 (.n_ena(w572), .a(w380), .x(w154) );
	dmg_notif0 g583 (.n_ena(w572), .a(w275), .x(w276) );
	dmg_notif0 g584 (.n_ena(w572), .a(w573), .x(w562) );
	dmg_notif0 g585 (.n_ena(w572), .a(w125), .x(w126) );
	dmg_notif0 g586 (.n_ena(w572), .a(w576), .x(w135) );
	dmg_notif0 g587 (.n_ena(w572), .a(w963), .x(w270) );
	dmg_notif0 g588 (.n_ena(w572), .a(w640), .x(w49) );
	dmg_notif0 g589 (.n_ena(w572), .a(w47), .x(w48) );
	dmg_notif0 g590 (.n_ena(w572), .a(w641), .x(w60) );
	dmg_notif0 g591 (.n_ena(w572), .a(w47), .x(w65) );
	dmg_notif0 g592 (.n_ena(w57), .a(w536), .x(w248) );
	dmg_notif0 g593 (.n_ena(w57), .a(w87), .x(w68) );
	dmg_notif0 g594 (.n_ena(w57), .a(w873), .x(w339) );
	dmg_notif0 g595 (.n_ena(w67), .a(w66), .x(w12) );
	dmg_notif0 g596 (.n_ena(w259), .a(w967), .x(w68) );
	dmg_notif0 g597 (.n_ena(w259), .a(w966), .x(w13) );
	dmg_notif0 g598 (.n_ena(w67), .a(w289), .x(w248) );
	dmg_notif0 g599 (.n_ena(w67), .a(w748), .x(w339) );
	dmg_notif0 g600 (.n_ena(w475), .a(w850), .x(w339) );
	dmg_notif0 g601 (.n_ena(w158), .a(w425), .x(w12) );
	dmg_notif0 g602 (.n_ena(w67), .a(w427), .x(w79) );
	dmg_notif0 g603 (.n_ena(w158), .a(w90), .x(w91) );
	dmg_notif0 g604 (.n_ena(w158), .a(w543), .x(w248) );
	dmg_notif0 g605 (.n_ena(w158), .a(w508), .x(w13) );
	dmg_notif0 g606 (.n_ena(w158), .a(w430), .x(w339) );
	dmg_notif0 g607 (.n_ena(w475), .a(w476), .x(w68) );
	dmg_notif0 g608 (.n_ena(w475), .a(w544), .x(w248) );
	dmg_notif0 g609 (.n_ena(w475), .a(w479), .x(w52) );
	dmg_notif0 g610 (.n_ena(w450), .a(w451), .x(w12) );
	dmg_notif0 g611 (.n_ena(w158), .a(w490), .x(w68) );
	dmg_notif0 g612 (.n_ena(w158), .a(w282), .x(w79) );
	dmg_notif0 g613 (.n_ena(w370), .a(w369), .x(w91) );
	dmg_notif0 g614 (.n_ena(w370), .a(w884), .x(w339) );
	dmg_notif0 g615 (.n_ena(w370), .a(w806), .x(w79) );
	dmg_notif0 g616 (.n_ena(w370), .a(w813), .x(w68) );
	dmg_notif0 g617 (.n_ena(w370), .a(w371), .x(w248) );
	dmg_notif0 g618 (.n_ena(w370), .a(w642), .x(w12) );
	dmg_latchnq_comp g619 (.n_ena(w93), .d(w79), .ena(w92), .q(w798), .nq(w797) );
	dmg_latchnq_comp g620 (.n_ena(w93), .d(w339), .ena(w92), .q(w432), .nq(w431) );
	dmg_latchnq_comp g621 (.n_ena(w93), .d(w248), .ena(w92), .q(w388), .nq(w889) );
	dmg_latchnq_comp g622 (.n_ena(w93), .d(w52), .ena(w92), .q(w99), .nq(w100) );
	dmg_latchnq_comp g623 (.n_ena(w93), .d(w68), .ena(w92), .q(w800), .nq(w94) );
	dmg_latchnq_comp g624 (.n_ena(w93), .d(w12), .ena(w92), .q(w882), .nq(w883) );
	dmg_latchnq_comp g625 (.n_ena(w108), .d(w12), .ena(w728), .q(w452), .nq(w451) );
	dmg_latchnq_comp g626 (.n_ena(w69), .d(w12), .ena(w70), .q(w827), .nq(w828) );
	dmg_latchnq_comp g627 (.n_ena(w69), .d(w68), .ena(w70), .q(w830), .nq(w829) );
	dmg_latchnq_comp g628 (.n_ena(w69), .d(w248), .ena(w70), .q(w831), .nq(w824) );
	dmg_latchnq_comp g629 (.n_ena(w69), .d(w339), .ena(w70), .q(w347), .nq(w340) );
	dmg_latchnq_comp g630 (.n_ena(w69), .d(w79), .ena(w70), .q(w349), .nq(w348) );
	dmg_latchnq_comp g631 (.n_ena(w69), .d(w52), .ena(w70), .q(w356), .nq(w357) );
	dmg_latchnq_comp g632 (.n_ena(w69), .d(w91), .ena(w70), .q(w950), .nq(w951) );
	dmg_latchnq_comp g633 (.n_ena(w69), .d(w13), .ena(w70), .q(w343), .nq(w342) );
	dmg_latchr_comp g634 (.n_ena(w88), .d(w79), .ena(w811), .nres(w249), .q(w805), .nq(w806) );
	dmg_latchr_comp g635 (.n_ena(w88), .d(w12), .ena(w811), .nres(w249), .q(w643), .nq(w642) );
	dmg_latchr_comp g636 (.n_ena(w88), .d(w91), .ena(w811), .nres(w249), .q(w368), .nq(w369) );
	dmg_latchr_comp g637 (.n_ena(w293), .d(w79), .ena(w410), .nres(w249), .q(w281), .nq(w282) );
	dmg_latchr_comp g638 (.n_ena(w293), .d(w12), .ena(w410), .nres(w249), .q(w413), .nq(w425) );
	dmg_latchr_comp g639 (.n_ena(w293), .d(w91), .ena(w410), .nres(w249), .q(w89), .nq(w90) );
	dmg_latchr_comp g640 (.n_ena(w293), .d(w68), .ena(w410), .nres(w249), .q(w491), .nq(w490) );
	dmg_latchr_comp g641 (.n_ena(w293), .d(w248), .ena(w410), .nres(w249), .q(w542), .nq(w543) );
	dmg_latchr_comp g642 (.n_ena(w293), .d(w339), .ena(w410), .nres(w249), .q(w541), .nq(w430) );
	dmg_latchr_comp g643 (.n_ena(w293), .d(w13), .ena(w410), .nres(w249), .q(w250), .nq(w508) );
	dmg_latchr_comp g644 (.n_ena(w609), .d(w339), .ena(w608), .nres(w246), .q(w774), .nq(w850) );
	dmg_latchr_comp g645 (.n_ena(w609), .d(w68), .ena(w608), .nres(w246), .q(w477), .nq(w476) );
	dmg_latchr_comp g646 (.n_ena(w609), .d(w52), .ena(w608), .nres(w246), .q(w478), .nq(w479) );
	dmg_latchr_comp g647 (.n_ena(w609), .d(w248), .ena(w608), .nres(w246), .q(w545), .nq(w544) );
	dmg_latchr_comp g648 (.n_ena(w71), .d(w79), .ena(w247), .nres(w246), .q(w607), .nq(w427) );
	dmg_latchr_comp g649 (.n_ena(w85), .d(w248), .ena(w535), .nres(w138), .q(w641), .nq(w536) );
	dmg_latchr_comp g650 (.n_ena(w85), .d(w68), .ena(w535), .nres(w138), .q(w207), .nq(w87) );
	dmg_latchr_comp g651 (.n_ena(w85), .d(w339), .ena(w535), .nres(w138), .q(w538), .nq(w873) );
	dmg_latchr_comp g652 (.n_ena(w83), .d(w79), .ena(w84), .nres(w82), .q(w149) );
	dmg_latchr_comp g653 (.n_ena(w85), .d(w91), .ena(w535), .nres(w138), .q(w55), .nq(w56) );
	dmg_latchr_comp g654 (.n_ena(w85), .d(w52), .ena(w535), .nres(w138), .q(w54), .nq(w53) );
	dmg_latchr_comp g655 (.n_ena(w85), .d(w12), .ena(w535), .nres(w138), .q(w822), .nq(w973) );
	dmg_latchr_comp g656 (.n_ena(w85), .d(w79), .ena(w535), .nres(w138), .q(w81), .nq(w80) );
	dmg_latchr_comp g657 (.n_ena(w85), .d(w13), .ena(w535), .nres(w138), .q(w139), .nq(w86) );
	dmg_latchr_comp g658 (.n_ena(w71), .d(w12), .ena(w247), .nres(w246), .q(w849), .nq(w66) );
	dmg_latchr_comp g659 (.n_ena(w71), .d(w339), .ena(w247), .nres(w246), .q(w872), .nq(w748) );
	dmg_latchr_comp g660 (.n_ena(w71), .d(w248), .ena(w247), .nres(w246), .q(w604), .nq(w289) );
	dmg_latchr_comp g661 (.n_ena(w71), .d(w68), .ena(w247), .nres(w246), .q(w600), .nq(w601) );
	dmg_latchr_comp g662 (.n_ena(w71), .d(w52), .ena(w247), .nres(w246), .q(w603), .nq(w602) );
	dmg_latchr_comp g663 (.n_ena(w71), .d(w13), .ena(w247), .nres(w246), .q(w745), .nq(w746) );
	dmg_latchr_comp g664 (.n_ena(w71), .d(w91), .ena(w247), .nres(w246), .q(w245), .nq(w747) );
	dmg_latchr_comp g665 (.n_ena(w293), .d(w52), .ena(w410), .nres(w249), .q(w253), .nq(w157) );
	dmg_latchr_comp g666 (.n_ena(w88), .d(w52), .ena(w811), .nres(w249), .q(w886), .nq(w885) );
	dmg_latchr_comp g667 (.n_ena(w88), .d(w339), .ena(w811), .nres(w249), .q(w957), .nq(w884) );
	dmg_latchr_comp g668 (.n_ena(w88), .d(w13), .ena(w811), .nres(w249), .q(w516), .nq(w515) );
	dmg_latchr_comp g669 (.n_ena(w88), .d(w248), .ena(w811), .nres(w249), .q(w372), .nq(w371) );
	dmg_latchr_comp g670 (.n_ena(w88), .d(w68), .ena(w811), .nres(w249), .q(w807), .nq(w813) );
	dmg_latchnq_comp g671 (.n_ena(w93), .d(w13), .ena(w92), .q(w857), .nq(w856) );
	dmg_latchnq_comp g672 (.n_ena(w93), .d(w91), .ena(w92), .q(w97), .nq(w96) );
	dmg_latchnq_comp g673 (.n_ena(w108), .d(w52), .ena(w728), .q(w102), .nq(w101) );
	dmg_latchnq_comp g674 (.n_ena(w108), .d(w68), .ena(w728), .q(w732), .nq(w729) );
	dmg_latchnq_comp g675 (.n_ena(w108), .d(w79), .ena(w728), .q(w731), .nq(w730) );
	dmg_latchnq_comp g676 (.n_ena(w108), .d(w339), .ena(w728), .q(w487), .nq(w488) );
	dmg_latchnq_comp g677 (.n_ena(w108), .d(w248), .ena(w728), .q(w481), .nq(w480) );
	dmg_latchnq_comp g678 (.n_ena(w108), .d(w91), .ena(w728), .q(w486), .nq(w449) );
	dmg_latchnq_comp g679 (.n_ena(w108), .d(w13), .ena(w728), .q(w106), .nq(w107) );
	dmg_nand g680 (.a(w936), .b(w187), .x(w782) );
	dmg_nand g681 (.a(w944), .b(w194), .x(w772) );
	dmg_and g682 (.a(w316), .b(w230), .x(w656) );
	dmg_and g683 (.a(w458), .b(w211), .x(w209) );
	dmg_and g684 (.a(w459), .b(w460), .x(w662) );
	dmg_and g685 (.a(w59), .b(w870), .x(w855) );
	dmg_and g686 (.a(w152), .b(w870), .x(w801) );
	dmg_and g687 (.a(w457), .b(w211), .x(w210) );
	dmg_and g688 (.a(w147), .b(w630), .x(w629) );
	dmg_and g689 (.a(w803), .b(w804), .x(w7) );
	dmg_and g690 (.a(w241), .b(w203), .x(w202) );
	dmg_and g691 (.a(w522), .b(w203), .x(w689) );
	dmg_and g692 (.a(w59), .b(w233), .x(w232) );
	dmg_and g693 (.a(w206), .b(w683), .x(w775) );
	dmg_and g694 (.a(w664), .b(w296), .x(w436) );
	dmg_and g695 (.a(w295), .b(w296), .x(w437) );
	dmg_and g696 (.a(w152), .b(w233), .x(w597) );
	dmg_and g697 (.a(w374), .b(w373), .x(w893) );
	dmg_and g698 (.a(w496), .b(w206), .x(w651) );
	dmg_and g699 (.a(w520), .b(w44), .x(w896) );
	dmg_and g700 (.a(w751), .b(w139), .x(w664) );
	dmg_and g701 (.a(w184), .b(w185), .x(w530) );
	dmg_and g702 (.a(w205), .b(w123), .x(w578) );
	dmg_and g703 (.a(w210), .b(w145), .x(w512) );
	dmg_and g704 (.a(w144), .b(w145), .x(w583) );
	dmg_and g705 (.a(w153), .b(w123), .x(w122) );
	dmg_and g706 (.a(w59), .b(w533), .x(w914) );
	dmg_and g707 (.a(w617), .b(w618), .x(w496) );
	dmg_and g708 (.a(w493), .b(w171), .x(w519) );
	dmg_and g709 (.a(w205), .b(w225), .x(w224) );
	dmg_and g710 (.a(w152), .b(w533), .x(w534) );
	dmg_and g711 (.a(w59), .b(w261), .x(w260) );
	dmg_and g712 (.a(w292), .b(w59), .x(w58) );
	dmg_and g713 (.a(w152), .b(w160), .x(w294) );
	dmg_and g714 (.a(w59), .b(w160), .x(w159) );
	dmg_and g715 (.a(w152), .b(w646), .x(w109) );
	dmg_and g716 (.a(w59), .b(w646), .x(w647) );
	dmg_and g717 (.a(w292), .b(w152), .x(w84) );
	dmg_and g718 (.a(w59), .b(w73), .x(w920) );
	dmg_and g719 (.a(w845), .b(w367), .x(w613) );
	dmg_and g720 (.a(w493), .b(w517), .x(w845) );
	dmg_and g721 (.a(w808), .b(w547), .x(w374) );
	dmg_and g722 (.a(w225), .b(w239), .x(w338) );
	dmg_and g723 (.a(w817), .b(w152), .x(w151) );
	dmg_and g724 (.a(w152), .b(w73), .x(w72) );
	dmg_and g725 (.a(w280), .b(w77), .x(w953) );
	dmg_and g726 (.a(w59), .b(w840), .x(w955) );
	dmg_and g727 (.a(w152), .b(w840), .x(w839) );
	dmg_and g728 (.a(w822), .b(w43), .x(w439) );
	dmg_and g729 (.a(w822), .b(w42), .x(w694) );
	dmg_xnor g730 (.b(w807), .a(w808), .x(w631) );
	dmg_xnor g731 (.b(w372), .a(w373), .x(w810) );
	dmg_xnor g732 (.b(w957), .a(w547), .x(w809) );
	dmg_xnor g733 (.b(w886), .a(w171), .x(w170) );
	dmg_xnor g734 (.b(w254), .a(w253), .x(w411) );
	dmg_xnor g735 (.b(w77), .a(w281), .x(w424) );
	dmg_xnor g736 (.b(w280), .a(w491), .x(w539) );
	dmg_xnor g737 (.b(w251), .a(w250), .x(w429) );
	dmg_xnor g738 (.b(w876), .a(w821), .x(w820) );
	dmg_xnor g739 (.b(w504), .a(w11), .x(w10) );
	dmg_xnor g740 (.b(w877), .a(w818), .x(w819) );
	dmg_xnor g741 (.b(w805), .a(w620), .x(w621) );
	dmg_xnor g742 (.b(w643), .a(w517), .x(w941) );
	dmg_xnor g743 (.b(w516), .a(w493), .x(w887) );
	dmg_xnor g744 (.b(w368), .a(w367), .x(w169) );
	dmg_xnor g745 (.b(w284), .a(w413), .x(w428) );
	dmg_xnor g746 (.b(w244), .a(w89), .x(w412) );
	dmg_xnor g747 (.b(w172), .a(w542), .x(w743) );
	dmg_xnor g748 (.b(w359), .a(w541), .x(w742) );
	dmg_nand3 g749 (.a(w460), .b(w461), .c(w221), .x(w220) );
	dmg_nand3 g750 (.a(w854), .b(w143), .c(w465), .x(w318) );
	dmg_nand3 g751 (.a(w228), .b(w229), .c(w241), .x(w240) );
	dmg_nand3 g752 (.a(w876), .b(w877), .c(w504), .x(w503) );
	dmg_nand3 g753 (.a(w128), .b(w127), .c(w569), .x(w568) );
	dmg_nand3 g754 (.a(w538), .b(w537), .c(w148), .x(w334) );
	dmg_not g755 (.a(w484), .x(w709) );
	dmg_and3 g756 (.a(w393), .b(w391), .c(w390), .x(w1) );
	dmg_and3 g757 (.a(w393), .b(w394), .c(w390), .x(w98) );
	dmg_and3 g758 (.a(w392), .b(w394), .c(w390), .x(w26) );
	dmg_and3 g759 (.a(w392), .b(w391), .c(w390), .x(w389) );
	dmg_and3 g760 (.a(w111), .b(w455), .c(w104), .x(w453) );
	dmg_and3 g761 (.a(w110), .b(w454), .c(w104), .x(w103) );
	dmg_and3 g762 (.a(w111), .b(w454), .c(w104), .x(w482) );
	dmg_and3 g763 (.a(w110), .b(w455), .c(w104), .x(w105) );
	dmg_and3 g764 (.a(w498), .b(w499), .c(w908), .x(w897) );
	dmg_and3 g765 (.a(w352), .b(w351), .c(w345), .x(w350) );
	dmg_and3 g766 (.a(w354), .b(w351), .c(w345), .x(w355) );
	dmg_and3 g767 (.a(w352), .b(w353), .c(w345), .x(w346) );
	dmg_and3 g768 (.a(w354), .b(w353), .c(w345), .x(w344) );
	dmg_nor g769 (.a(w694), .b(w439), .x(w438) );
	dmg_nor g770 (.a(w416), .b(w406), .x(w405) );
	dmg_nor g771 (.a(w407), .b(w406), .x(w256) );
	dmg_nor g772 (.a(w529), .b(w528), .x(w649) );
	dmg_nor g773 (.a(w629), .b(w177), .x(w178) );
	dmg_nor g774 (.a(w503), .b(w624), .x(w625) );
	dmg_nor g775 (.a(w663), .b(w891), .x(w167) );
	dmg_nor g776 (.a(w571), .b(w230), .x(w237) );
	dmg_nor g777 (.a(w558), .b(w207), .x(w208) );
	dmg_nor g778 (.a(w909), .b(w900), .x(w899) );
	dmg_nor g779 (.a(w844), .b(w644), .x(w495) );
	dmg_nor g780 (.a(w287), .b(w288), .x(w361) );
	dmg_nor g781 (.a(w366), .b(w230), .x(w238) );
	dmg_nor g782 (.a(w230), .b(w175), .x(w231) );
	dmg_nor g783 (.a(w522), .b(w241), .x(w648) );
	dmg_nand7 g784 (.a(w699), .b(w702), .c(w697), .d(w928), .e(w397), .f(w788), .g(w401), .x(w400) );
	dmg_nand7 g785 (.a(w699), .b(w698), .c(w697), .d(w398), .e(w397), .f(w402), .g(w401), .x(w696) );
	dmg_nand7 g786 (.a(w706), .b(w698), .c(w701), .d(w398), .e(w700), .f(w402), .g(w401), .x(w399) );
	dmg_nand7 g787 (.a(w699), .b(w698), .c(w697), .d(w398), .e(w700), .f(w788), .g(w789), .x(w695) );
	dmg_nand5 g788 (.a(w267), .b(w266), .c(w264), .d(w263), .e(w235), .x(w567) );
	dmg_nand5 g789 (.a(w267), .b(w266), .c(w264), .d(w793), .e(w235), .x(w268) );
	dmg_nand5 g790 (.a(w267), .b(w266), .c(w563), .d(w793), .e(w162), .x(w841) );
	dmg_nand5 g791 (.a(w267), .b(w266), .c(w563), .d(w263), .e(w235), .x(w262) );
	dmg_nand5 g792 (.a(w267), .b(w265), .c(w264), .d(w793), .e(w162), .x(w792) );
	dmg_nand5 g793 (.a(w267), .b(w266), .c(w264), .d(w793), .e(w162), .x(w161) );
	dmg_nand5 g794 (.a(w267), .b(w266), .c(w563), .d(w793), .e(w235), .x(w919) );
	dmg_nand5 g795 (.a(w267), .b(w265), .c(w563), .d(w793), .e(w235), .x(w234) );
	dmg_nand5 g796 (.a(w267), .b(w265), .c(w264), .d(w793), .e(w235), .x(w842) );
	dmg_nand5 g797 (.a(w267), .b(w265), .c(w563), .d(w263), .e(w235), .x(w913) );
	dmg_nand5 g798 (.a(w267), .b(w265), .c(w264), .d(w263), .e(w235), .x(w645) );
	dmg_nand5 g799 (.a(w493), .b(w517), .c(w367), .d(w547), .e(w620), .x(w619) );
	dmg_nand5 g800 (.a(w267), .b(w265), .c(w563), .d(w793), .e(w162), .x(w163) );
	dmg_nand5 g801 (.a(w632), .b(w631), .c(w809), .d(w810), .e(w621), .x(w622) );
	dmg_nand5 g802 (.a(w744), .b(w429), .c(w428), .d(w412), .e(w411), .x(w958) );
	dmg_nand5 g803 (.a(w538), .b(w539), .c(w742), .d(w743), .e(w424), .x(w423) );
	dmg_aon2222 g804 (.a0(w731), .a1(w482), .b0(w487), .b1(w453), .c0(w102), .c1(w103), .d0(w452), .d1(w105), .x(w937) );
	dmg_aon2222 g805 (.a0(w482), .a1(w481), .b0(w453), .b1(w732), .c0(w103), .c1(w486), .d0(w105), .d1(w106), .x(w767) );
	dmg_aon2222 g806 (.a0(w350), .a1(w831), .b0(w346), .b1(w830), .c0(w355), .c1(w950), .d0(w344), .d1(w343), .x(w768) );
	dmg_aon2222 g807 (.a0(w349), .a1(w350), .b0(w347), .b1(w346), .c0(w356), .c1(w355), .d0(w827), .d1(w344), .x(w939) );
	dmg_aon2222 g808 (.a0(w26), .a1(w388), .b0(w389), .b1(w800), .c0(w98), .c1(w97), .d0(w1), .d1(w857), .x(w781) );
	dmg_aon2222 g809 (.a0(w798), .a1(w26), .b0(w432), .b1(w389), .c0(w99), .c1(w98), .d0(w882), .d1(w1), .x(w2) );
	dmg_aon2222 g810 (.a0(w545), .a1(w546), .b0(w774), .b1(w775), .c0(w477), .c1(w175), .d0(w478), .d1(w651), .x(w650) );
	dmg_or3 g811 (.a(w36), .b(w38), .c(w716), .x(w717) );
	dmg_or3 g812 (.a(w36), .b(w37), .c(w25), .x(w440) );
	dmg_or3 g813 (.a(w36), .b(w442), .c(w23), .x(w22) );
	dmg_or3 g814 (.a(w767), .b(w768), .c(w781), .x(w525) );
	dmg_or3 g815 (.a(w937), .b(w939), .c(w2), .x(w3) );
	dmg_or3 g816 (.a(w36), .b(w778), .c(w779), .x(w433) );
	dmg_or3 g817 (.a(w426), .b(w644), .c(w649), .x(w610) );
	dmg_or3 g818 (.a(w899), .b(w898), .c(w181), .x(w144) );
	dmg_or3 g819 (.a(w36), .b(w40), .c(w192), .x(w193) );
	dmg_or3 g820 (.a(w36), .b(w39), .c(w190), .x(w707) );
	dmg_not3 g821 (.a(w528), .x(w527) );
	dmg_not3 g822 (.a(w420), .x(w419) );
	dmg_not3 g823 (.a(w417), .x(w418) );
	dmg_not3 g824 (.a(w416), .x(w776) );
	dmg_not3 g825 (.a(w6), .x(w5) );
	dmg_not3 g826 (.a(w206), .x(w378) );
	dmg_not3 g827 (.a(w376), .x(w377) );
	dmg_not g828 (.a(w232), .x(w475) );
	dmg_or g829 (.a(w644), .b(w615), .x(w614) );
	dmg_or g830 (.a(w896), .b(w7), .x(w6) );
	dmg_or g831 (.a(w626), .b(w9), .x(w44) );
	dmg_or g832 (.a(w239), .b(w240), .x(w290) );
	dmg_or g833 (.a(w175), .b(w176), .x(w633) );
	dmg_or g834 (.a(w246), .b(w598), .x(w737) );
	dmg_or g835 (.a(w648), .b(w594), .x(w593) );
	dmg_or g836 (.a(w140), .b(w139), .x(w295) );
	dmg_nor g837 (.a(w291), .b(w181), .x(w182) );
	dmg_nand5 g838 (.a(w623), .b(w887), .c(w941), .d(w169), .e(w170), .x(w942) );
	dmg_xor g839 (.a(w244), .b(w245), .x(w612) );
	dmg_xor g840 (.a(w517), .b(w493), .x(w971) );
	dmg_xor g841 (.a(w620), .b(w893), .x(w892) );
	dmg_xor g842 (.a(w547), .b(w808), .x(w894) );
	dmg_xor g843 (.a(w373), .b(w374), .x(w871) );
	dmg_xor g844 (.a(w367), .b(w845), .x(w825) );
	dmg_xor g845 (.a(w284), .b(w849), .x(w414) );
	dmg_xor g846 (.a(w280), .b(w600), .x(w740) );
	dmg_xor g847 (.a(w172), .b(w604), .x(w605) );
	dmg_xor g848 (.a(w359), .b(w872), .x(w741) );
	dmg_xor g849 (.a(w77), .b(w607), .x(w606) );
	dmg_xor g850 (.a(w254), .b(w603), .x(w611) );
	dmg_xor g851 (.a(w251), .b(w745), .x(w415) );
	dmg_xor g852 (.a(w956), .b(w692), .x(w417) );
	dmg_or g853 (.a(w666), .b(w416), .x(w858) );
	dmg_notif1 g854 (.ena(w232), .a(w231), .x(w13) );
	dmg_notif1 g855 (.ena(w209), .a(w558), .x(w48) );
	dmg_notif1 g856 (.ena(w209), .a(w46), .x(w562) );
	dmg_notif1 g857 (.ena(w209), .a(w765), .x(w135) );
	dmg_notif1 g858 (.ena(w209), .a(w851), .x(w126) );
	dmg_notif1 g859 (.ena(w232), .a(w773), .x(w91) );
	dmg_notif1 g860 (.ena(w209), .a(w762), .x(w49) );
	dmg_notif1 g861 (.ena(w209), .a(w761), .x(w60) );
	dmg_notif1 g862 (.ena(w209), .a(w561), .x(w270) );
	dmg_notif1 g863 (.ena(w209), .a(w592), .x(w513) );
	dmg_notif1 g864 (.ena(w209), .a(w208), .x(w65) );
	dmg_notif1 g865 (.ena(w232), .a(w238), .x(w12) );
	dmg_xor g866 (.a(w171), .b(w613), .x(w518) );
	dmg_const g867 (.q0(w14), .q1(w47) );
	dmg_not4 g868 (.a(w897), .x(w626) );
	dmg_not4 g869 (.a(w862), .x(w509) );
	dmg_nor_latch g870 (.s(w749), .r(w633), .q(w632) );
	dmg_nor_latch g871 (.s(w867), .r(w663), .q(w499) );
	dmg_nor_latch g872 (.s(w532), .r(w334), .q(w147) );
	dmg_nor_latch g873 (.s(w150), .r(w151), .q(w75) );
	dmg_nor_latch g874 (.s(w614), .r(w529), .nq(w230) );
	dmg_nor_latch g875 (.s(w519), .r(w614), .q(w520) );
	dmg_nand_latch g876 (.nr(w656), .ns(w143), .q(w759) );
	dmg_nand_latch g877 (.nr(w182), .ns(w816), .q(w183) );
	dmg_or3 g878 (.a(w36), .b(w41), .c(w473), .x(w693) );
	dmg_or3 g879 (.a(w36), .b(w42), .c(w43), .x(w31) );
	dmg_nor g880 (.a(w8), .b(w144), .x(w501) );
	dmg_nor_latch g881 (.s(w8), .r(w7), .q(w9) );
	dmg_dffr_comp g882 (.nr1(w47), .nr2(w47), .d(w309), .ck(w311), .cck(w312), .q(w46) );
	dmg_dffr_comp g883 (.nr1(w47), .nr2(w47), .d(w121), .ck(w311), .cck(w312), .q(w561) );
	dmg_dffr_comp g884 (.nr1(w47), .nr2(w47), .d(w120), .ck(w311), .cck(w312), .q(w558) );
	dmg_dffr_comp g885 (.nr1(w47), .nr2(w47), .d(w550), .ck(w311), .cck(w312), .q(w761) );
	dmg_dffr_comp g886 (.nr1(w47), .nr2(w47), .d(w217), .ck(w311), .cck(w312), .q(w765) );
	dmg_dffr_comp g887 (.nr1(w47), .nr2(w47), .d(w216), .ck(w311), .cck(w312), .q(w851) );
	dmg_dffr_comp g888 (.nr1(w47), .nr2(w47), .d(w549), .ck(w311), .cck(w312), .q(w762) );
	dmg_dffr_comp g889 (.nr1(w47), .nr2(w47), .d(w330), .ck(w311), .cck(w312), .q(w592) );
	dmg_mux g890 (.sel(w122), .d1(w330), .d0(w120), .q(w308) );
	dmg_mux g891 (.sel(w122), .d1(w120), .d0(w330), .q(w879) );
	dmg_mux g892 (.sel(w122), .d1(w550), .d0(w549), .q(w766) );
	dmg_mux g893 (.sel(w122), .d1(w549), .d0(w550), .q(w447) );
	dmg_mux g894 (.sel(w122), .d1(w309), .d0(w121), .q(w456) );
	dmg_mux g895 (.sel(w122), .d1(w121), .d0(w309), .q(w866) );
	dmg_mux g896 (.sel(w122), .d1(w217), .d0(w216), .q(w485) );
	dmg_mux g897 (.sel(w122), .d1(w216), .d0(w217), .q(w445) );
	dmg_nor3 g898 (.a(w529), .b(w891), .c(w144), .x(w143) );
	dmg_nor3 g899 (.a(w663), .b(w466), .c(w467), .x(w460) );
	dmg_nor3 g900 (.a(w530), .b(w531), .c(w844), .x(w816) );
	dmg_nor3 g901 (.a(w616), .b(w496), .c(w655), .x(w908) );
	dmg_nor3 g902 (.a(w178), .b(w179), .c(w176), .x(w177) );
	dmg_nor3 g903 (.a(w594), .b(w522), .c(w226), .x(w225) );
	dmg_nor3 g904 (.a(w861), .b(w594), .c(w204), .x(w203) );
	dmg_nor3 g905 (.a(w438), .b(w437), .c(w436), .x(w435) );
	dmg_nor_latch g906 (.s(w546), .r(w737), .nq(w773) );
	dmg_nand4 g907 (.a(w695), .b(w696), .c(w400), .d(w399), .x(w929) );
	dmg_and4 g908 (.a(w706), .b(w702), .c(w701), .d(w401), .x(w727) );
	dmg_nor3 g909 (.a(w134), .b(w133), .c(w570), .x(w569) );
	dmg_and4 g910 (.a(w77), .b(w280), .c(w254), .d(w251), .x(w540) );
	dmg_nor8 g911 (.a(w77), .b(w280), .c(w254), .d(w251), .e(w284), .f(w244), .g(w359), .h(w172), .x(w422) );
	dmg_and4 g912 (.a(w616), .b(w654), .c(w166), .d(w165), .x(w869) );
	dmg_nand4 g913 (.a(w230), .b(w500), .c(w868), .d(w179), .x(w180) );
	dmg_nor4 g914 (.a(w611), .b(w612), .c(w414), .d(w415), .x(w972) );
	dmg_nor4 g915 (.a(w606), .b(w605), .c(w741), .d(w740), .x(w739) );
	dmg_nand4 g916 (.a(w9), .b(w10), .c(w819), .d(w820), .x(w506) );
endmodule // PPU1